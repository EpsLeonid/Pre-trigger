XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B�M'�āVmg�jF���f��O1d��.�oT�sk�鳗���V2���E�����7�S��;�� mxs�}w2�S�X��&d�X�6A:��3�U<�JV��=nu<��(k�ݽ��|� <*��c>œ���ј�l�ؕ[��/'&��rcN��8�d$���_ݖt���h�~Gȍ܁�S`�^)��QB�}�����f�pVi�Ps�xh4 W榪�5L���w����A���;����$@���Ν����'���iS,��0�p�E�����k8}cq���$0�~��}�Kaθm
O�T��X�7��@�3q߮n+rP�� ���5���O�A��3B�<�t�n�*�T�/��1�Gf���9G�F�+�e ��J5��l�]NG�k,I��E���Y"q���"��^�l9�oFW�(
e_G�?��F-m^ ��&n:��!�!.C��� ��Fb�i}CC1Kd�x��[���m��	���	i�?�럼���Y�O����ͭ�g��t>�V���.�Ǉ+h�$7�:��W<6�%�������-��(�6؇5i��qe��l��zS~(��H͉}����39'�+S�	2����]�Mm�n�#0^f���oYCiNܝ1��B�)-E���nU�,T���~RveI�J��1�A�j�	��\3����?�/�n�3|nb//2m���߷� e��U<^wh`Ob�B1���9k�h	qhHi�IZ�K��2"��I=[�<zđ�v�k�C�9�XlxVHYEB    4071     db0u=	�H���� �;@ ի+�V�kr����0Z�w��
.�Ҕ�����P����K���/:����&��.�X���+:�@ܰ�>G�D��7m|�nojb!���Ύ��j�#�Gd�N�=����Ǩ"O�V�y5s77�#8_��v)0�E)n�<W�y�Lv�)S��s�:�`4֡��F荇t֖tĝ�_HuB�O�{�b(��I�`���5ݩ#�$$��Jsؑ��B�"�/r�mdu� C�/v����ڕ��y|��;'
Z�>UR�A�oE�W`3(~ݯ�bM+�&n�/g�Φ����:Y���|UÕ�����G��V�h��V��\������-���b<�;��<i���^%�����Զ�E�Ry���/�@	����)�CJ<f���FK���J�޴F�y6J�(qh��^깞|(����PɄ�Κ>�-C�����ߟ���3{�vQlK�z5Z�X��m���T�_�t�ُ!�z��gBݢ�g���K�Il����_��B5�`��^a�E�䮅�U������Y��Ú*��w-"�����"v<Ğ��G�]V&;ȑ�)�����r�w�{�.r3�>���,D�OUN��~T<Қ۩T�ܭ�=�
��r���,����.�l7{' �+�7�]S�������V�0ot#��a�|G6OCj>�@xk>?Ϡ��(B�5T��]�-H�>����7r)���㆚��ԑԵ��5�Z���K7���u�rg�R�q�0����8�9���� ����E��T�կ%��,4 �c��g]dR@���붢醾�l��AY%\[�h�8��|q'e�@9F�������Q���w:QZӨ)5��wB�,~c�������~{]� �8�xqog�Y�z��Y�$*ܽ�;A^E|����\��j#����]���;��O=f3#3��:�|�����+�f7���g���Յ(�u�~IkX��U�g	��/�wu�Ge7 '�]X{��B���Ǟ~��� ��ޣ��U#�BcO�	�C�-���~�wo���~$|�5�YT0n)~21�o��W���%��'�gB��=$1D�ʓղEhr��":��,o6�ɑ&f0���z�ٰuaOH�У�;6y.�����ηm�ZQ>�Q#ދ�w;'Ĕ7O��q>僻-'��Gq�5��Vqp��F) 	K��O����i��~�f���j�4A-�<m�#�ՠ����L��x]��k
�<v��K���R�'���Kiz�Oˬ�2�J�ԪQs�Rc�6��s��QQs���ʪ���&���CYR6@wp�������@�h�"����!)?��s������q���X�N6�*C)��c����2��P����ד�u,��v��'\�s@OE0�j�L4�����H��#��'�B�pb�(�sL-�)���L�5���jNf=���Q�����>�����l�� ��9��ԓfb��b���s��b�H����@��v�CV@��,rS����>���FIu�w[߷�%hh��ӵ*k,y|�}F`'Pe(��~��me5c-�-^���F"�	�'����KM	���!�ӆ�BD5�s3��87�Q( �;u�F�<
ߞ���C(����̐��^ݞd��jp�=�l��7Q�n�еR
�C��
�F��3��۵�j�|݌��vB/�R�������� &�L�%ܸ+�	aEݩ���Ch$��K�� 4�tΨ��s�M��<3��=Ĵҩ�|�ݾ �Q�^a�H�'/CJ��BK��C�%�ښ|��\X'� �1+� Q�w�Ì�g,Xl�eiwrOu��ܳ3[<��TQM3G.UL^q~%Ź?
_�^��Y]�ɥl�'D4=�zL��U��-��y�,��|E�+�'g����6=�����j�<��Cn�B�j�`e^TP��o�p&�ETBY�c��
�
5��*;�[G�ԅRG�i��A��^nU ���52�D����6a�H��7�H�#ɨ�m�h���� �p�B7r���Ef�!:h�~a���K,�����K�����P���"2lZ ���<�����A��l��4���8L4JE��-�dvjBȅcB#F�*��e�77���!���Ύj.��������p�8��`>��#	�Ed�Z!dֶ��%�Lb����棍x ��$v���~uR�EY :�1g������FÈ��$����쒂��b�F
�4�Y>�ϧ���'E�v�h���?.�tDo��TSeڿ)`7�Fl�m	6���X�hx?��-�b9NQ�R�K��S��Og��&L��jG��_A�z�+�g���l	%F� /���*h������Z��u\���+Q_3�q��[�� 
�-�=���x����K4��%�0e`L�S)5>ꝶ;oYtL�H+�5�n
4�~�'�\�;U2�иJ�%�$���Â�v���;��� S�V�ϭ�x���(�N1��?8�#/��j��Aʸ0�/n��d�)��<>�d��#8�KX��o�����$T{haф����1�LI�\�[�h�2�!	�ى[�Mo}����k�Y�9zo���t��%]�, �Y��`���f?�`a���A�?ʉwE�c�f?�n�Ɠ}�i�ab <�8�}7��j�y����X��d��d9��b��>m��g����IL�����R>��B�Hk�6L%��bT9����Mވ�#>����7���<����D6� "��ό��0����!_\��Y>�y~�y�1��!��Ȑ-''�L���k����	���3��	��hd�9�0^�q��غkq��a	���Kd|_v�K��Ί~��v�ոg[���n9�
���0�A��۩��oxW/� LcS��	��īȀ[��c��c����_�6�ߋ����bX�G2��N��o6TB��`cM�n��i���9SLh�^RW٭��s#�������'�j�>�==md�mH?<f�DD�.4��i��d���j!I��ڱ��y����J����_D�HM�H��Pdū�S����ΐ\����3^��-�X��oX&��T��(��.��t�q�wP��ܷ$��˓P�O�˨���ݶD�7?޴�` ��T�*�o���gl~���d�*�z���}��yC!#���*��-Y��I+w��Κ�{��]��Q�n�����b;�HL�j���
n$�w�ܹ

>�^�oXB`�7�"^>q`�bsc�꜅G}��+)�8������;���Hn�N>�t��,#�]��u��U@�ǖ�faE)U8R[�Q�ÄI]H�\�ƥ�������w��7B�$��	W�L,� %�o��<�_4��E0��9o?����T���&�]Z�EY����N� �	�iu�
����阮l�'ˈ��B!Q:�n%��5��he� d��I&:�D�V�)Q�~h'�c����Ya�aZv&���9a\I�