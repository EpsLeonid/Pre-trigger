XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��J~4%'F$Q���uN�o�;Ŷ�n@��ޗLyJ���>*dԠ`7,�(�ރn�����G�$�%��VW*m`b�o!��mL�)+��r�M:�q��g�2���B���D�q�*��"���]g[��d2�m��/�Bl���\أ��cc���8J��@��S��ۉ�7�¹�PK�=���,��nb8��iH"��Р��x_j=R�N���*��p(э�=��j�,|S�q�&35��w��C9�]�$A��󥆩3���v5�Z����pZ��� -G+�� �1q�߹P��� a�c�����nn<^�F�4U�bJc�>7�c��ZU<8��Z>c�BY�����\��)ڗ߬O�Ѩ.����i:\@�ssʈ��[r�O��pj���?)�c�k>���l �{N
�J��"\E�6�1h���yV-�w`[?�VoD&!���}{L����[��46 ;�骒�YnB����*>�J>�X>�6�p�)�ZGa����B�����b����hJ$8���Y����[~姗G������s�φ?�.�F�_.�9#/��{,�*��d���3�K��=CRA���4; �/]�/� ĥ����n6��� ɦش.��皵@�ơx��4il᭗�|S�v�{lL�3����K��f���ѯ
���?�졵|�yؑLv�1��.]���c�Y�}�{uh�),KJt��I�;0T�n��@[&5$�y���S0z0�E��l�d奠x���I����-s�7�XlxVHYEB    38a4     d00L?�ۥ%//�)��F����? ��Cn����:�k>����8�%1�#�,G�����b�'V��z7sT/k�6�����o�w���3v��&�}d56�]�:P���J��83�9�#IBv�2�q�*-X� �Աoz
�Q�x�aO�QB��ɗ-��fu��%��f��U��QE�`����[-�fZ"��A��DW��]��uF5`�T����1"����8�Qza7�x�tҤ��ݺHe��Yuڌ��d��2
�3�qGz��]�Z�C��
r�\��<¡���z����2�ߑ\ӕ߫Q|��m[抳�.xYOX�6s��5�$r�y��Cۉ���<Ι�JA#�@g8��j�A�.Ih���T��a���Yx6hv<08�,l�����y/nK����;��������g��Kť��.Ո6!.`�� ���5��j?��AR; ���Lm^a�A�A
��b���S�Zj(�~A!�����SU��#@�0�ꏶw��e3XJ��4uUZ�偧��Hv�����ʍ�P��U��`��!���o?�E;�2��2\�a�̔�ή�ĥ*�+q�dQ��rZlNdª`	�e�.�}�-�2e�+�w�M���Z�N��>�����7�-ҦS|����tx[�ζ�`(��e�!k18d�kօç�qQ`��n����,��U,�|��:^�K��0��i�E}���+q����� �|tY�T��!��@Ke1�'5�U[�)D1n��I��v4:#�_�Z�I� �40Q-�N�߬|�͑*^�����(��]����෌� �-%�S��2�u7h_��l�=�B����ԣ-k^S��ڱ�ki�|��yD�^ԺxW�S)�ߘ�D٘^���k�,F�a�,.�|h��BD�u%q�/\�Q�-�vC�`��4��]�p�����g�����!?�X���b'+#�/$�h���/�ֶ/N_�INp��wlh�u,	�#��;� �6��冯#�b0L ?�$��������;�It�.���/����\�t�1!oo�K�#��zh\���1�sCj6�����Vy�myhR'ۉQ_�80i�
v�@�I���^f>s		�|��WMf��������!�+8Ux���9�g��j�1����O�u[|	19킟*�y� <�)��mh�i�[�ww�fc"Ql|-��h�SY[89]5�1��Y������� �D�����f��ː�M8.����1�U��M��,�:�Y�z���F��:��oSDn�G��	H��3�W^�ҡ�k�D�Ap�W�vA(1;�G增m��g�xZ�<YP1�Ȝ������$��Q~����0'�XJb&c�}��'���Mm�����d�`�jt�T���ֲ ���X�S�
i�ϥ�T�㎧���2INM�k)���� ���j'��l:A�2a?4�ޫ��B��b���f���<��0�\;Rv���b�I����Uȯ%~gc��7{u?^���y���v�R2���/0��Z5�g9)�[N�T���-h��G@"�sFz�1��gp��_:"����à��A&�������������=Fc��]�]����0t�"-�ܠ�T���w%�/p���3�9��4��� �Z ���w5G.��^|�?�����G�5�Y?�Q#-|���{�y6s �=�T>)T�]��8�I��;9EZ��)nH����
Q�y���s!:܋,�>M�x�Ve���e?x2���qZP硙ޖ��"7GM4=ŀ�ۙE��5Xh(Tc�ΐ�vŻ����)����*U��#�Ӥ`��6���mj�n����h�-# U�K��1t��,=*�D��� OB��m]��^��=�/��i��,��S��_lĚ#v�Ɲ$���{�k�%N(�`qy��n�A���# �5�_����w[6ޓ��o%fc>��>a�?�9_,����2A���ۙ��p�d����6:�����_7���}�
�b���f*��Ю�.�LQSw�f�wrY�=���Ї��Ǧ_Q��;��U��$[,�e[�\6��7yL�g��5��2���t����(*Z_�� 8�`�@�����x��G�)�Kw����y��c��6G4� �L���=�Y���(8��)QK�M.ޣD�+w!P���ߦ�%�#c�F�>���_ ߖ5�DJ!�= �P���TR���! �\ �FF	1���aq�h��)u�;}��[b��܇���iS.�$:�I�Md4wm�!���њ�:�y3��;�M�Eښ&�U�mf&�tq�t���p��_��񼴼�M�:^��]I� g`|�S�m�Z9�^�ۅ��	K!g�¹��"�.	l�M�^�"��d������H��A��i���Vyw�Z�1C\�� �j~D�����Ě#�קE�b��ˎo�<?�w@�9E�R�7�edÔϤ��^��x8b��Ǥc�������C� I� 2�i�;��#uP��o]=��Y�,8��/
�Lq��/n$���~�wp`_5���V�I3���P����D�����d�p?��hLi�F���^k�����د:^-Ƭk�%�4���VK�(�a������ՕQ��˱8��#K��o��޻��Ï�yK8�����i�v���{[z�LRRp���5��N��ĥ*Q�����!����40�8Ǧe�=:��%�������i��dv#�kL���2�!�	�R>����J�ċ��
�0���o�"��oƞF�b	����2ֻ�h>N���rY���2���0g%n�RL�b:]�ʚ��ٷb�g4�\g:�*ζ�\�M�C�Q����}W��EY�YU��Z>t9��.E]H��a�guHL��sy�H�͊�Ƹo����ٌ��R��1�l����X��߭�^:���zΗ-B8C�;�6�
��V�Wu8�ƌ�}V�S�d�{B��$��]+�m u����%�� ��<d
F��S����n1rP!���G�vo�����ލ��s����܂�x!�'
����G�\�!�'>8��6Wu/)"H��d�<�;k`ȥtg���n�`��V=G�14V:�p��ŽΈ �P��˩����(
��T�����@[���.m��(^\���o��&���R�;i�f�y�#UAS��L��[rc�~�=�5��䂃����ڌ�N������Q�;��"����]�/� ��e�~�I����Xb'J��%��E��`bȼi�i�