XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z�O�Y��;�="/����,��:�(Yݖd��'�j��[ڑdr����y�Q�h>>`x����-ѳm�"Td�[׾�:�QJ������������O�,|�i�����[;�V�b5x�:37�&��f-{�v�n5�$ʹ���T�و�cW�;%��Z�-	H>/�$q5�YB5ǵ�4�à������^�M�*rb�X��h�����zy�<�������$�����/��TrU+]N�/w�<|)�L�3��i}�@��p��u��e���m�[����s�F-�|��d/�0�-gTC�(��Q*⊹��
����!��Z��@�� 5W�/�� ��ľ��Jύ>����$8{b���l��{�{}i�_�[Fy��\uU�, `�����`�C��z]F˶hCH�2������(b�m.$#T�����JG[
�k�
Ԯ��yL;Z����`*_�^�����W&4�H?�p�>�Bd�u�0rʥ��ӛƟ�5�,qˏ�&�2��D�T�ll�d������u��hkJ]�A��oܤ�a��n��i�Օ=���\'�@��&=fL���g��4��q���YWܖW��5y��-O���рE��Rp��+�5ވt-$���d����e�Zz�X��,NV���1B�/q(�l��1��a�/㒃���� _ޘC�$lD�k֋�k��@�7sH4V1X4��l�\V�d8M�,Jx�r��u�6\|Wc�l��ڛ�{L�R,�B��魿`*&�XlxVHYEB    4071     db0N2�7K�l���V��L��+����_2�RL�u"H�1#�:��"S�j�����K-����6�u�^o\JT�8�9.=��gY(���61ƛoa�1>N_OY�-J��O� �w
�����({>�pG�S�2/���%���C�J�ſ:o�C��J$;�C�Zwt�د�	�P�'K�怫���-O��h�)�aW��Ĕ�)��p:���3I�$qV�|)C�Q	�;��5dU�'W�;��E�B�X��y{�l�O� �f���U�i0��Зم����+�]d�A�l�@%Z�Z ��m����L� �$T�q4��Y��K0����`V�[��<��闬���Od�T6Cɯ+�.]f��s]���mVx��u��;�WZ
��#3�P'��{�qn��͍<��<h�X�~�۫6p�R�ƬJ��1�f6�5yeA��K�I�ۻR�y���f�ە�!z�{{e�*�q�5`Ҩ�mJ�������0Ls��=t��~m���|�� �u,��YP\����1���E��- t���書<"mY[wX�v����-����C�������!��@l�H��w�TN���ݙ�?Z���-����	��8v�J��u	�M�h$�-n�|��A����n:�C��Ә#��fnT ؑ��5�+�a�ԅ$���_XV�BA����(Kd?/9�k�����7�P�t���.5ź���d�4G�
���$}R�����բ����O��t� ,���F��N8%�]b%B��IaD�š��M�m�U�٨�+_ņ����i�U��4�����OM��*ve%(���.��b��!T㒖��j��g�.��G EcV��T
E̜A����?�z��F��AE�xO�,M�p��17	<fz�v	�.JF&�⡓M�э=l8�s�d�G���8Ô9���'�_�c�.��KB<�ǹI�nF>o���I/�S�}I10�?�>-�S��nF�d�g=��a��0{�:����h��F�{f`���:�e��h�V�{*�r�|��bn�N���"��VarB_��A�q���SM��a�rR 	���gǂ��b���d� ���CW��~L�΀1)h���|p�8���-�B��_�p�"]�ԣ��ѐ틅+�ՀI��dK4�'���z!Ϟl�{�����>m��[�`F�b{E�.����݌L�x��0z���X&���U�&��T߸:��FnE�R��gG3s��Z��:�\-�4�-,'3�b=��/ث����e���hB����ˤ��k����YU��4���tK�2���}G�)��lu:gFү��O�m���r�EI�l/Ҽ����ꡕ�8͈��O�Rn~��r̵<�yd���M(E��@�C�/��E7��������V-'Me�X�W�=�4�Z��+7����Z��acθ'�J�:u���x_J��2�:�ŷ��ħ^?�6�qAO�r�눙�H��Z�^�~�ًl����m��M^y�x+�Q^7g �;�� q*N��>��D�b��'���{3<��	��x��֓c�݃����i��#��-��L�>�=�/_�+�;
@��Yr���7�E)�^s�B}R�w��Px'p]o|��w�	H�]�xC�$�ZR�y�Â�~)��J!�M�[��"9��Ξa=��{�2b.���l'����d���f.��. !=&�E��:˂;�D�>w6E/�T$�+�4��i.�����rn}+�;�\�j �Թ��^�J^��>Rjgzn�j-K'���0�u�> �R����OKa �3~�iρ����aΝ�K���`X�vl�� ���^�ꯔ�F%�la�.�ew�L�l�u|�f(�Оѡ�m��7�������؋�i�M��*^�ŧ����
2ֿ�ǀY����;����3T5�C���;�Wd�l���|v��=b2�S����?�I"��B�����0#f���[ŻO��Adr�w0�v@�՛��F1D�,����3f�%o>f"�A<Ѷ��2yJ.�8"},�y���.�ܭHQ��z�x�߉*�|ۤzxo�t�l�qk� �����U��U~5�Ɛf�֠�+�@TiBx�q݁�G��.�ӡb��I<l��ՎIk�1`m/�n��x���E�@�i���4��r$d�v�W3C�7zO� MqG�M�kM�6eqNi�.l|�1Yѫ�X��ݳ�'�h��Wg�����av���E��&�V�� ����U�je`�l�=������e^#���i5#GK6{�Ġk�#�`�E�ئPw�c,g��˦O�O�8�M���y��ȈgK�_N-=��x�R���c(&��6�9��O+��/7�:�h�|2=����'ލ�kK|�������-��)2�E�{R��2���P�@�Vi��G�bbR=�ț-،�mo��6�`j��^�]r��"1���+�8n)y����=�>v q�������$�ҥ�a�t`y��6�H�M�}�L��㗆���jH-l���_4_�У��{�!P����_J��}G��o������?�V�.�9�	�R!;���j������$����@���F�Ҳ�̤���28���O���JF���M+�:��	��[�M?�BKT�s �Vw��� ]��ϴ��s�?����gZ�M��K���*��v \�W�e�X{E����)�1S��O�u
�LL��<�+�'.e8$�����᧛�)i��{x~��-���xYԘ�k�$�9j�x��Ko�.��V(���)s�ښ�����eb���6D��2���V˚�Z����y��CQλO
����ޯT��'���=L�IHM�Y�U$ �a�j2G�<Cfz�*�&,@DF�˫!�Ü<Aۮp[	ja���;��Ioc?��}����H������,{X$?�x��n���q�Hw�V6��Q �c�� 
vD����� 2wi�v�C��W�i�����fw4� G��o�šx �����ߙ� ��1��;ul��
��i[��ǱE��^����k�B�딗,8����*��{VӅ�������a+��[H�UX^�C��\r�Tz��S9pխ� C�lP3U� �!�k^Tb�� F;�v�BH��1`�Р�nJKL�����:Y(NWx���J[�z E�+��������ġ Phۨ�Xt8;���#���g��F�嘬Ǚxs{��j�L]3n�J�JYx�V��}U���)^o��.�ƞՏ�6�8�`�ļ�	NR��Q���J��\{>�L�Q��MȑclO��r��}���1(�`�M/�l���ѡ�W�[�aĥwuq�h}�bv$����7x�Aw�l�Թ�|9Dһ��G�5^"�>^ѣ��y=�`F{a��T�5����ru 	|��� jX���?]�v�(�G�[�b^��ۿy�ү��9I�51���^�Q��eΘ����}^��