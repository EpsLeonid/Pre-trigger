XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���M`%b�D�N�1�a��x9{a_��)m��O�$����A����\o:���/��ɴ�"���Yk"�����ۓ�$f������p�<
Ҫ�F�\*�_a����Et�,�`�I��/,o&�h�P���cShA몲�Zi�����7i���SԦ.�EV���fuA�N)�����X�����>/lLC��[�y:�ĵ9��s�ea��,�Dp=����m���xJk�Hz=e	�N���(X�!:�� %X�S��ٽog�x���4V��<�F(A�b$PX0�}ΞF����O��2Շo�>d[Cqm*�lѶ�j*l�*���������=EC�9�`�R��X���pW�xb��Ń����i��ȵ	a��e����&Č޸.��?������� ()���>ѵ�/�����t�h�IJ��.���@���J0���J��f�px�r�0��(Ԍ;�_�i� �@Qu��� ����p�|��q�敹M -����x����X����}�A�
��r&������=��b�e�@����L�{�O$�{w�5�I�~��%�e����V~��	��
t��Z$
u7�iu(�x��� �z������x-H�����| hm�L�����������%�~�|�9��3�D���.8/�G���庉78a�=�`�=�{IA_p2v���e��G�׎uF�m�B����Ag�%z���oy� ��nڽ�X:����I�pRZ\#��ї+�f/JȾ�l^XlxVHYEB    2fbd     d209������\�FD:�L��k�w�|��	
O2�e���|��g�"xZ�$�pOW�����+4Ѕ��UJΣ���X r7+�,���ʗ��*����;��p�3�ץ��E����٘�Jj����<TiL~c�΄��L��#�hL鏑�D��`���JȂ�4��/e���}�ҟ�8bT��-ef�d�� �/����r��3B�Aܵ]�y��9*���� o����ǭ����|i�p�&�_aT����7������١�E.����B��N��������e�[�뼦g�>jI�f�t�I{���O��K��=/�^�#���<�SB��@T�	�{�(ؤ��N|�X�lr���#1![��"��YL���k�K�k��P�>�..;����Or�\�O��[d�$]ol��b�&V��C�vi��@KLc����¶�]١(1s��	h�p<�i=�� �9��z�}��V�'�ВYw��N�"yBc.}/wO�͸9��X@Y\����������7���Q(Bט��3�c�q.R6�/٭���7��Z��gB�*p>���h���ֱ#��N���h�,��i[�М	���<�2�y�,x�و��0Mn���Ƽ��G����N���Gev�]��=��rdL������!t 8~I�����)����Q�HW}�Hܖ�[�C��I���R<��l0���m�]iq�lQB$�9��8�;�C2;������@����y�^�.a�\��l�5Zv�Ū�`��-=��Jm��G�}s��fG��_�J��c�{Mb�����~�W��t5X��T��C�3��/Oއ����'(C>$�s\
nK�pbsy��2?�9�A軙:$�P"���{�4��j"�/�H׽��҅��"ћk"h���C�P�n�AǸ;<��G���f=v�WS�f�c��$��Wָ���s�r$%�O�X_L�Wv�=5�)�asBQH1��}����4Py���T�}{ٝu~O�9�>�����Rffi���������0�H밽�M֮@{ܸ7X��E\��q_'2���4s��-T���c�Lļ~�±Us��	)�G�b�v�%��`�̤o`4O�U᠎,6�!�ʻ� q��t-��n�<^�Y���������7�f�����'V,��G��ף��{�&�Ą�?fs�&�JQy���%�@͌��J�Q���羴JÊ�m�cS6'� �j��A��dɇx����SڄKE��(��b��~aJa��"K��*�g�f�ۡ��hI�^�ȏ��T�8�����2�N���5���;P����p�>|��IE�;W^i��x�覜�F,�;���R�E�O���CC�O`d���ٻ�ˀu<q|$�����#_E�v����I��R�o}Qu���"��K�n=�;�Ώ�?lr�͡�g]���`��7-7����Y���T=�.p��AuPW�P�e����.�Fz[Y������;���3�}��[RW0
�;
��U*9����	���"	�z�$��=��4����^���IRK)2�"�[gP����d�}�;�B�Lf��g����w��l���G���t�P�yc@7g���~rs���6��=�Z)ǎ��_��g#$z��6�=gn�4�x]W��>5��42ʑ�����^x�oP��fFG�!�U1��9'3�ɑ��	`[6��m-9s�s��{��Ow`PU�SѤ"G�2[�{���F��� �x'��H@ʹ���n%?IMzx6p�/s&���w�t��g۫a�o/?}���:ϨWI5��Z1r�%kT�h�En�݊~Fp��i��_�� �؋:K;���7��1��",H?��>s��)�6:�-QN�X�
n� gd>!�1�n�����w2^t�,�������',�v)bu��03;�e8���ؓ%��1�G�ߍ%0������Jc�b����.�㕫��[��Ĝq��ח���d�8�|N����0j�d��=�+�[,��ܝ`�P����K[�C�^X;/�J�4���g�3K���ː�������j}#�xGLG$Fw��׳�)��(p�Ē��e������5a�'�����M�Q�4n��9�<�F�����WB�<� x��p=�4U�4���Y�/�a�8����8}�N͢Wy�q��Ш`����|(� ���ɭ�\��Sa�]�.��{����l|�鲱��&���������k@��&c��$�8�Sv�L"x�����n����ɇ̎�}\N�0HX�+Uy+Qn��Y��.t��2�S�KȌ��l*D7�ߚ��� �k��婎�

��f����~8 L�ׅ�B<?2A���\���x8��It%�0V��5�=�B�����=��F�91q-�PPUVX��l�ln=��L�]�+�h����ʖ�y����֮z�/x�/(���~���C���*}����[*�ڭd:q�8���s<�K
܁��?�J������斊�����7�w1���F�2�6T�d�ϒN|�f̔����$
pF��R����B�p�C��/�l�%�8#���#�B����s�˟Ոkv��`�'*�%���F�E�:�nޥ��|8Θi��űs���X�����#����]�ҷ�"��R�om� (O����q|�q�|��U���4,�L�D���of���� ^O�<����;� o�O���ͺ����^ 8�Œ�~UZ�8��2E�տY��*Ty}�Ө�B|�^@�$�
k��ٕ�V,��g�-k�BF�j��S?�U������
%���"����հa�}�z�d�d٥��M�2�'�dV�r�Ҭ����x�j��9�^Rχ�=�G5����M�"(h_���@*���b%��R2~;"%pB��6�St�&�&��501Xѳf���BB���9�p!$�&&��a�ȺUc||�2d�9��'�e�K?fa���]a+�c�A5\e/ ���`�	�x���0�׳�2>�{B�A���7n�+CB�]����.����+�	!� Z�03�,Ob��j�|���4FOl��M�WYt��#hc��ձ�Z������7���I�Y>=�lx�D��J�L�fb�M���;�$!!��5¬By<�S$T�墫�#�E�2��V�4�.��(���FHS� �f��=�2���#����"m6��QƬ'���o暋=�9l�-<���|�,��2�Q3G����V������k�|r��	��
���L4F�aQ�&���h���0-!{���;:�(܃�