XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������\~wGnI��ST�^<%���K��ϕ�Pq�m��L�Q�m������5�S��7�W\AAv��m�=��R�} ��5R�lb�yމFM2��ŉ	�{o�]����xfC��8���n341a��x�O���@N`�k%��r��|�S�:�,1/G�^gڊsuW�<���x�tZca�� ��{rk=xZ��P�&�?	E���� �ɉ��R̋Hg}�Z�[O�I�����`���V0L��N���1��Q>��݀�<Kd����g��U�4[��r(H��?�ٍ��q�Й��j���"�k.��kNEf��0���
�w�,�M�����rR�[��e[���f(��?аR"�fyl��z���@;O�e�BD�͢K7\�9�M�a;��b�s�`�	r��m��_~���$S���Z^��|��o����ߡ��d�
<��h������e8����j/��A�Y�䆿"�������)1YE���ֵ#��U�͢N�M'�`��%�ʮ��Y�_f{M�>���c��������� �W�lL~2F,T������������}?Ǐ����<$r��Ws�j���G���-�~�g�^�*'��p�A��J���@��>�����YH��9
fz��p�������`Ǹ^&��"��ti��TĶ��k����`d��ްJ%��] �S0�L�${9G���:WL��7����';ʱd�4��/��*�EƸ��d�A"�pK����}��v�:x��]�l�iXlxVHYEB     f8b     650��Ƒ��wN�U:8?� ��䨍���ǀ�E.gZpJ@��"�OP)�^b(��Ѭ�Js�5��h@S�%u|��v,3�@2���U~ ���w�$d������R���"�"��͎G��N�*�8�M*��p�Vz R�d�E	�z;�� x���Y$���Z�g@�ʇ	�n�%�T�t�رR/�e�Q�c��%�)M0b�:R�w���I�{�M��%�W����A�kA�.I���V@� ����)��!�mQ9d���g1�h�8�=���˖���z�~�&}�T��6���3.�'���"r������IQ#R43�������g3���a�'�0�ڼo��0BWc6d�f�z�w��NYy�8!�l��[�� H�lH��I�)�ߒK:}	���z��9�������	��_^y'����x�s�.��k�+�t�� �8Ki��浘�h4���Q�l��/�9��پ��-Hg��P�c�V?�L��5�f`<	-�9�<���\���i�^�����>��sʛ��Eg׃<��2d>O�L���ZK��Nar]h��|�^ܨr�T���P�e�Q��Uuhͫ�P����ėӴЊPL������
�Azv�VI|�Oh�^�c�~~j?�U�	�/BUV<.��Ԋ0�͗$�&���C��&k0�ϋ.@q��U�� ^?9�Y������#f���]�>���X��S���&l�N��+l�մ��K�jr�rw!�jf�����\�0�N����x
ۆ�u�G��^�^�m������U����:��f�N��k-��r�O�UG.���w�iU�"0˟��Ds������֌@w���W�\���=�H���If�v��H���ض%�	N�|���bb�	�R��[���u�^=v�jf$�M�Y�?�����^Jρ��B��Yd`�������,\R�߱���\8jҠ3#��ݓ�����6[���7�?]�<��J���c����Xd�9[.�����������hR3@(5�r.��LSW�s�Et��1���l����d܁E��N���U��{�e�ڪW�K}à�]\d*9%#��WvǳR�4.�Q�ڦv'��Z���n�<��Dn?���'8^��%s����e��(%+Û��7�T���U����ڲ�8R[v9o��~6}�� ��W����S�o��K���MS�D��OȀ���5e���骱�G���6Cz� Fshx-f�	^�z��FE��/�H^���׽��6WdM����`�z`���V�6U|��
��zt�v]"~˯�6�,�܀��xꙏW�9\@��\��"&�Fv�]����ӷF�[�a�&�l�F(�7�5e��G�D3�Xe��)�����86mz������(�o��3��e�熘������
��ӷ�-i���H3�I0�w�>RNI�q�NY�"�E����B4����Ђ��L({q@��(����\�I"���i��׊�a�O�"i� �^w1�}](`�:�U�#�� a��;�AW�K��}�s��ՃT��@�~d~�����.�A�v�|������HT ���@Лˡ��b�