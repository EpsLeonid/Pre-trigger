XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���[�� P�"�L���K볞`赒z���e�!l���A��{z����2R[3$��G_��?AH����퓕���M�Pt���#�WD� j^����
���0nEi��Y��$�!7����2�^���VI�S>~�@�A,������_HŖ��D�wӇ9�@�HY�����>���7�fj��e/����;y����8$��W��^��'1G���vWK����!��4+*x�>���Mi���Yu�v��E���5���/Z�:����L���@(_OՋhW�+����IG#�!����|����S����c����#�ݏjg� �y�^gd�ّ"���pH��E�'ҼV��kn�3dOJ��$��w�a�Ai2*��gM#�FMK�vg�mD�@���^�t�hD!m W|:��������H���m����e5�V)��Rqe�N���kWp*)M�]Jgv�������5�d<�CUi�M��q�\ە�(rcQ��QV��$���	W�7O���	ۥ+� ���R���"5��MVx5�_�Q��P��P�(� !󣊙Ǽ�&ꤡp�E�3�d9����T�X�w�+��3��uDL�#n�l,��E'����p j!�i(��h~�>٦r�n���يrk1�Q�-9M���Ku���n��DB&�E�#7~�/�~��!SVIy7�d3m�$����j�!7�(�Wy"tV�4Kd��K�A9(o>Bj���̜�Sd7�lS�hJ��LXlxVHYEB    159e     7e0;��:��3���?KL�����ɽ�	c*8"ۜ7$�r���P�z�xv�����9v]�El����}����#��*�2V�S[Uy@�R��ֹ�M���|o��Z��S�����:t�pv����0��7����NȂG���R<����6g�R��L�q��*���'D&�At <.���&����-5����)��M�{p&�z��pn8��bl5�1>3X>��c�l��d�=a)��i�>m�t����w{b�b�>'����i�e��ʚh�t�k郮���WR��E Hvl�H�/ ��>񁻠��_g'z��h���{��_��sY�����@nJ�TMTs�T�P�Q�<�����?�ľg->�}b�h�̾��.<����WwsDD�ⰽ��M͂'���Cp�ϱm�̲4��]/�c�ҽE&Ic㇤5+��T��l�-� ]^F�� ��F;��82~(8�u;T���ٗ�Q%(Y�M��3�8�˙}za䢥��`-Jf��D|�6[�*s��K�/�nTi[�Z8Զ��
|k@�@��[���^7T
E����&�
���I\DiK�;pa�ⴕ+��w܁0��˗�d��,)=n�u��N�O� r�>O�a25t�nD��H��X�b��\,����)�\��L�Ѵ��[l�k�)�y
6B�J�������jK��:e���#~:�3@ے~�d��V"r���2�CF5�'"+��v�
���XԌ���@o�Ο�R��E�@z7�m�|N9����uVU����O%���ѥ�W~�
~p̸�E��R����;���qb��3i��q�]���)!�v���lL֜�z�XP\�d�����
%����׈O��W?�$n6Ki][K�����'%v�ǑV�4�eŐ�����p�O�ΉٹN��8����ud�6º�n��m
�Lr��~~�E����m�-B9��σu���8�,Ҋ�J�Q�0�=͠���;�/Ig"���(��t��4������Ob��@�WĬyZš�9��j5w�� �qh%rc�Gz�]�9�Wzt=Қ�-e�P�u	Uh�̅����Ot� �Wq��Cb�/Y ��N���x%�]��B���n[Oi�gnrYהGHz)Е���M��k��%y�G��b�f(�:b����YLLx8ӹH�J;ɽ�D��q����ui'e(�Z[)��[-=�v$ݔO1UE�V٥���'���'�⡙��m�Qsú�j�%��㑫p�'�F��l�4�[��g�D���
����<���Vp�yo3�O�.<��=��q�g�G��2UОL.�r��Ps�r����ń�뭑��6��yZ����_�\��~w@*�ƒwih��� �"z���Nt�n'ձCk��G���Ӣ��?Z��%�Ⱦs�#AxF��T��J�7j�+������:)V�}����%q��f����oa9$�
TwK_�@�a��
d7�v?$l�2��I��� �J��D���d�To����_���Q@n����!��&FC��g��!z+?���7�3!\����ƶ;q [���-��9<�w�m=<��M��Y?^D9FVɽ�ǁV���S*�����굘�imΟ�xK�[����U'6
$�Ю� ���%!ټn}���0���a�.O�'�G�";^�Ͱ:9��qV槿��&w�q��ۉ�];1ޔ��k,7�gK��	����H[M�l�}�V�QHQ����;<��Ð���p������g�����AI`�VS-������;	g\��p�����y�'�}��K���}�U��_�\�/��y��5ׁ��9FV.x�b�n���G���L�vV�P�eY~(t��`̰fPzn7~�x���hG��d���|� :$��i^��6�lڱn��C���!'L}g��﹨[7��uI٩L��da