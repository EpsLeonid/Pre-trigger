XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Mv$�d]P��	��W��V��x�-JE��)�`��_�	ܴ����w�2(i\S̷���Tq�8p��T$}�_�2��[����0��n^v�eR��V;��\�g��8�{t�A����]s��?�Vt�aO�ìC\��Q!��ɹ�@�/��:�����Ψ]��+m��0rSĺ���^�1)�hs���%lN��l�Y��0Q�I��h���3��=�~���E{�NQ���yd�2J	E��.BAV�1��M�z%� �-��������,v[I72Y�I�@��Dz
U�s�l+��po��ѭ+�9p�7�G3z�!O$Q�,�$p�g]#/��WƮMf~m�&CN[����{� �m���BP�����5Ņ�R��N@�\3�f����6sLw��$���mOq=��?V���NG��#]��aFSdCWH�F,i�h�%�IJ�D7F�OӪ(�h�~x޹N�<D��mVbl��������L�����]�q�x��x��`�99~ՠkn+K���4�z$��}д�L� ��s���& �!�O�C ��weY����o][�S��d�$ve�x�j ��W���p����x���?�܎�i��	B
M�6�u�J��8|:���Q��������/{�|�+
�(E.?i����.�B &�HO�n��R7��E�٬e1��Љ��u���o�GJ-G��6��{G|���l�Ru�5��[���a��!��h^?�3����^�_X��XlxVHYEB    5571    1410�	�P!��P�od'�8߄0�^�"7�Э)9v��#B��׵tQ���'ͯA��`�bBȳ��+�7>��B�غ�*�i��/.HV�=���\M�3����w�N�8�� �Ɉ=?�fU#r��R����,b|��Ҽ�'{a���xD�UՂ��6�|4���b���%�^5���b5��ӧ[��µ���	�.���O@&�$np$�]��b�g�4Lɠ���n���H�z�Ά����Ý}���Ü��GS"���@ZD�mO�����2w�����I��u�J�+z(����?Vy|>v0k�<MF�lS5f�W�,���͚����3+W`T�rh��gB��ۮ:��HF�;�k���+)D��v9�H�pYT�a%�[!F��U�[�dK���+�SUŹ	�yL1������ ��Cǳ$vv�i����
��)Dib�?G�?A͊�m��(��sr� ��W����4A��\q�;����Հw�u^t1�c�;�P/�ɒ�t��NaX�zG[�" X�T0�:z�"�6��N�~�P�k��v)��^������_%��f�]�~�.&�5l^M���DC����;��W�>��c~�˛����Cҵ	�(�	 Mzi��]���!��B磔?^E,=Q��Q�o���d{���~��+���I�=4@kͺ�|�b4n���:��_~D��ޣ ��Ғk򉮅�ecq@��_��v������0(�U���:�؉&B�^4���? e�ϭ��9�oh���2��A�<��V���o? �0 j4��C��� J23�#R�E�����Np�b�z��f���+s	��RY���m4���k�B&�n_!xo$�G0��ɨ��@�y�\ډ�
�ʢ�M?��7��n@�3������W�yΐ�K�%9��
3��i���	1�m�t�Be��1C����l�L�	�ٯ%�y$�D�#�G"!�4L�FV�@�6µ�~�{6���?�Ć��)�{��O$[�h����x��rg������j����%K�S,iPG:lKO������i��T?�/�au�\DZ� �\�HĹҢ4v��YQP�N �vJF#�L��t4g��K���J�e�{�U|����NW�	�A�%@�;��D������?p���X�	�aN�l��X�*&�]��(9(ŷ����!	�C��s��6a(�Ц���j��u��F6�c0Nz�c�:�/�������pu�+%:Ӳ2g����n� n���N��	%�_9��v��H��K�^~䩎|8��o��Ld�/@̫mm+�B�2��+YJ,xL�,Rz9�臨W����}��K7�3_X�D=Z`3��T;!0���
�Քy� ��-���8�]��	ѝc�B��F�!���-2��H\T�
�JC���oI���%�?�����b�����Xb���)�$��~)����G������bEm�������"�x�wK8�4j�YX���ܷl3l�XFd���4� �������(�;R)GE�sW���~[F:�n��=d�M�_d0�v�T����L<$(&n\���?���"�7��4t�u��)��xѴ�tn�a��3ᕃ�@/Q��#�b@a�"��&���ᐨ<yG������5�<�D͆[�+ۭ{t��e �m�Wqa�~�~�w�-���W�C���}hE�T>��?��C<6-~�>�cG��㗗�u�T{Rq�DW�A�������{��'~�{�)��/�|G.��gv�wz����I�D�[��vQLA�L�B�
+��U.́�$���)�͵
'��6_A�J�����PެM�]�=��'��R�����s`��|��F_��� �e?��;֥V�F7/klRp�����)+d�4��u�����h�e(��ˏ]�=T��\�(�VD)v�yl�R�ȶ@�u㏴���q�l��N�]ɏ�����	�3J���a�JqXEG;�6��/'�{�Ӱֶsz�����[�p5#���ŗ��Ǻ��)DM^A^��kԐ�Lst�N^4���

��H�Θ-H���p��y�@P��gp�WηR3���*.����|V�	2���s�/�\��Z�d?BG㢾 ��w�8�6l*;�:x�]k��n/7��ɻ�F0=����s瘮%�*�&S�3)RӢP����~�dAW�䦒�=+�H��8�:=���<�j��g�~1�K��1E��{��_+�}��=�o�т0zT����)p�e��U��R��(1���
)3���� ��ʥ�$���n2����1����:a�\q{:�/V2�Ҿ&͸F�P��a<�!�dNl2I>��P�;��u���Ol�s�����
�Eg?ofb!�����<�1�ۤ������A�.�c��m@�=/�|k5[!�v��D:�\�(�}�#/Uh�<�CA�i�U��\�FD�+G���%�5�b��Oik�����S��ڛL�dF�4�j+�J�Dz��1�~�إ�Ӟކ,l���Ùԙjta������|gy�-]��$?���-7!���
��w��b̋J:2��M-'o�W-,n�Q�m�]G��¯�8-NE,W	X(���00�]e;>q�`�0@��_
�VL'm�,M���t��sZ�Kr ]��[O�|9�yv��j��b�����u�?u��^@�U�����r6�ʶ��*߁<�;G�s� E���pUx��C�Ǹ�܂i0F�f�E0L�Cc�z��H>�xWx���;YCf��8�\��
�p�s;oYt!X�Ș$蝚���O(O�9�U�;�}gP��´��|( �%�Rob��5��,1�'��G�8�2���[��qs�6�3��9Oj��h��r��S�K뿦)���wF�+q�*J�B0A.��ˌ���]/����98�H���_a�u�x�<�b�k�r� ���P$�:���u=��h8짗��v"!40'1�d��^��yR�?���\O"~+@S�r�������W��[�a�b�_e݈��<3ra�d�ˇg]���J�؄*�hH�u~h�ѹOS:P9�ϕD���f����>	M��hK#zB湇��>-aV
�
">��H�񖪯�UI0���`������p�Xe�ײh�ԅg�20�O��¢NJ���y��Ob��(T6O�,�R_�7�Q�y����N�����6Ӆ�HH�uK��\�~"U��3������I#U�]��O��yts��vs�6��m�j"�ڋb<���ɉ��t���� �_^xis ��S`��G��#��tå�y���,OU	iK��cߤb�6<b��+f��ʗ=Noq-mY�7�73%[zSVI�e!^K�*�j^?�4�CV���R��le���d)�,Z�+�k$;���$�R{
,X �n��X�c��z�К�f~���[���t�E�+�������H��Cb����~G��m���븷�<�`hl�r���Ø�*H-^X;��j�0��� �(,n���y�HP�	�"�n;�1�u�sP��}����|���%�;�D�^C̆��2e�[lS����aKM�3R�r��@�2*��J(���P��Y8��	��~�	,צ-�WI�NUב�X���QL9�^-R��+>u��/�Z����*����!\���Ǐ�T4���B,�;��p�b�ٌ6���-�R��o�u7jC�`G<k=�I�
М�+�yͩH#S���xF�WM�uZ�:�W>D�1@΃������+�X3����a����;64"R����-+�ˏ�NQ���Xb�N*�8v{�ӽ� %&��r�'-	ĀGD��%��ùT2��Nw��(��Sb�%������Q�%��N����+Rq�͹j�=��
�AF�d���n�oX�0�9-�g~��&��ⲷ��E*gfZ�|���)-��.�{��M����[^��.�~43-����HR�܃{��k�Ұ'&��V�e1JK��B����M�\�p��g|� ��&#)vl���2���a*Ec�����~B���Js��Q��@΋����3�D?����,��*܊�&_�5�Y<6䋮Sz�s$Ϙq���)>u5�C�C�M�+�ã��!����0�9��F�z��+���$�[�̦k�z�^�0�D���2\>��'�qC��g�^$��䂫^~g����2�j�@(b\;�������G�rY<�7��x����Hd2�����B}�����	m�o$33(�lkf�ʄX���ٽ�W*`�e*mF��츛�_�O�s&����M6���R���V$1C�*\������w҃���,0���~>Φ
{�8�\d��ㄡ(�MW��.�)e' ��������}x��'���3���� �j���t�$�jK}f��⨤�|H������|ME����a�.�y ���"���5 �j%�=Ph}�����h���Q7���7Uy\L� ��{z(�K�ϩl{�C�\`�!�w�͎B+�����<Su����g�OeE�dv&�A��I%/-��oe�=>�#6��.��aR`8TD�1�V�d����	-�L|� 0󭺽�WR~fG�t��a�s�gE�<Kz�#"ԇ~U�Np+-EFx&{:�Uz�ҡ��|L�� �,�e5:��q��5W��JPU/y�V� �4����,~X3��egG��U��p�دw'�o�XN��~���L������j�oj\fR���ӑ{�x���ZZo:<����,��#,��1�k�����Kr��h$8>�w�^�y��?.�ˋ��vt�G�8mo��oNĀtfdQO=����"Ti�y�C4?��2�gf�o"B%��av<�������{@��t6%�W���aa���/I00��U�B���v�6�&9md,[a	�w%���g#y��G�7�Ԭ�Hn~.?������w�6����yS���?��~���Z��/�l����A��' ��b�����PMt���_jg��"�)���%����we$:k���K��u]}�||���@�@�T��:��4�|��Q#�����