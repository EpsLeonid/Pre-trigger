XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����J�"6`�2Q�iq9�!�kLs �8M�ԋ_�W� ����Z��$7s��j���"?E��)��<3���7N~Jbx�FH���u%H^x���
Ø�>��[���
�n[��R�q-���eK8v8Q;p��K����㽶�{���>�堺v���s��7h�%�BѤ]�]*�y��~ў��X�Vn��4yB=-�3ۧ�.5�D��Q'GML��kh��/��h:�/�$�Ն�灳����:R���A�n��Q��F�.#2�ظ"� Y�n1,r
W�SL���!I
�!IؚT2�qC���D��%��*�MÅS}y{�,��,2I�
Mq�j����i,�!��1��\rY����Wj�T�w�ↀ�$E!Rx�"�R�?C����ɶ3f/��h.�R�6��>:��>�������޻�l�c0%�o?z�ތ϶��nh�4y(����?4�P7�Tx���~�AF���UE9�{�t�3m8~�_����G|
�6c@Go&�A���gmL^X�t�/$�� 
��t�$��f"*�Z�jD_��GO(�κ�O6Y{�����N\"O:i��vZ���>�#��\{{
�f٫g)Y��>���F>R���ra�
t	�{>��u��"P����㡭%���́j���t�Ɍ�P�t^����i��ӸI�Y�jK*t�}i�c�����A�������\��lf!!%D��Mh��">ٰ��,�]%�7a���(���5a#�yl[�|p�j�1���f"XlxVHYEB    1a2b     8f0*ܞo�"R����~����m~���!��q�Ì���[���g8���J'�:y�����O���N.� I��wh�_���T�#l�\��ǩ<-�OH�?݋��\6�VP�%�.N�/���Ѓ�f.#
ׄ��a]�&�B��"��s���P���������i
�9r�^}&KNq0�.�DZ�o� ����������w]Ҵ�^����e�y��ϋ�IFe�6STT��a�M掊�a]!����,4���oK�O����N�����d8�3։<�4�HpG.����d��a���z�0���> D�.9vj�!hЪ���&�8DfE��r;�d�����am'6E����2�}0��`A�����ls�^;�r����M~%5嵕i�Q��U���`�茕ob�<�h+��K����65��u"���]ȿm@��!�7�H�Y�4�ٛ�����/?L�-S���Y�Xe�B���p������,&7��_e�P�V�B|k�VѿA1*��y����-]c"Y7���Q�SO�_�8�Pn�rbi�W����������2�#C˵�Ϙ�	�g���� �7��ϦT�ʹ�bD���T$L� YQ`�Ʌ�TP�6&cjk�y��c�}Y�1H��1U8�.}@'y6��4������&�=YpL2��s�\Su[P]6�V��L���쵬��]�/�8t�E�\�:���Fq�,`�m�5�*!���R�[�q�����e86k	"���ĊW��6.�EPޅE��A�?�߾�J7��ɑ�>.�(��k*��r�^/�B-�:,Ô��{I��E[!��LU����I|���/�4	ok0�dr>j�a�g�{�z�ԬCr�\�t��,�r�W����ϰ�l��GՄ�}�wV�`�Q|�����09*�*��rfR�C��oiO�5����m���g��B�ݳ}0�ʒ���r�ȉ�3��ٴ�^�g2�����$u�/
��gv������b����g<T���2�]?K��:���+��TF�#���O^��_;��-1P������6�uB#�U)_ ��Z|�{3�I]�F7���zF���n̊`u��A�t7=	�yz�B��T,���{�9�.��H�~�[�4y����[µeX���٪��i#�Zx���lm�W2�]L�ĝ��`���bi��$T-vϯ��������h�@�&5�!�4/�bQʐu�Kő�_�u�{�䳢��3��~Hm!�P���(��v��L�v�uL��.6U}��E9�@�;b�dn�Ӌ{�C�3}5���0���X�O`�3�d�(�uD�Y=y�Gs3t�dۨ)m�=^Ȓ�������#L��|u8fF��O��޼vo�^�����#|!��VZ��DR � ;fȬ��� ����k`���G��]r\T"ؚx�~}�zd�r����ۀd�8l�����Q_���-\���)"\�A�*��i6ژ�!S���X޽�X�ӝϺE�1�b�o� �A	����Z��;'d9j�켿�� ��pr�5�Q��" b���)��T��:%TP�]/�/���as��c�V���jf�U~�ڥ��s�*��QC��k�$^�K�r�������pm�F��y���R&(Fl|���f���FC�%���d���ޢ �40��5�pV	p�Ha�٤�'J&(J�^֣�D��M��h��𠕝%6v�N���!b� � �ܜ�v���@�(ڴ�R\wA�96��L"�fڮ�Bͩ�I�1���}�n�Yޢ�5`�N+:Ӆ�O]��tr  �ꯎ�:u��e�m=b
�=�F��mZճ��� �)�*�3����ܯ;R� �G���vvx,LD��wg#�홓��(1��`��w���b�柭����ܠAP%sN�k�����E����7Y�@����ʓ���g���a'7tbC�����m2�~B��+л�`�v���{f�Ê)�C�� �d�7��0�~�S��X ��@�sb���[��s�hp����Eq�"�kP&t���`�:O@��LN���R��{GӢ.O�m�Ϡ7e
6�?���B�|o����cSf���V��'��MC��~�7$$�鏔HJ;� ��uW����cYD��e�K'8��Bz�l�v\*������x��'�	�[���zF��
`���}�ڹ�G� �1�=�=�Ď��<�[����1)Q�����ia��&���̑�5up�������