XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^��& ���k�1�$����Q+�º�f'�\@*!uDqA@"'{��%X��EFٌ���WnЮ�a*�i�`�Zy@�O�E���:Pk����j�/����S�ăx�� O��M��[q�Z��S�}e~A��G�aNy!�`:�
K���4��U������hI�d��
����:�la/��Yl��`��������!�23j����8�h����R��s˧��k�K�^,���0�+_��f4t��Zi(	�;y�E�8s��V�-���%	X����1�]�N����Ͷ{v�t��[���nn�PuL[��3���SGJM^���R�|A���ʭ�re��:�C'=���l�!��{P��b���x���$c�C�	o��R�lAAX�֠#݌a��U��\<2a����*i��JO�7�k�_�
�+ԛHO��UӲ��U����F���o��tJ6�����-�6�*;6!>�ǭ�W`�gBIB:�Y�Ŭv��FK��_SF�jږ"�j���l�X1@��s���S�"'��"��M��{\Tq�H�=�A��At?s3��2>�YX��� �V���k?Q���Xܿ	~t1�&��{P����6��D:PS��27�������S��������<��)z�ED:���֝�
��W�ˈ���?�W���4�S�iu܈��p�h�EBt��θ&d�V�H��3�s�}#��Ca�9�R�	�=$�����*<�)nL0m�C�O!A�*,nB�a�XlxVHYEB    1001     6c0����K�#k'��N$NI�ʌ��u�d���1�D�&�V2�R+���_�U >g�tԜ|sSO��5l�˛�@��A49#s�CM� ������H��`���xס�y�	����'�l/�x!ʂ/P\n��Z��$�{YP�V�0��H�7k����-t?,�Ps�a�}�`����{U���))~�K�ﻅ��V�R�#�O�gQ�.51���˷�E��*Ҁ������~�UDo���1-�C�aU��-g�w�_K����*QC�V���k�pK�Ğ�1u�}���J��e+D��z���pѣ�)��D1P�Om�>`e�1��h�I�H=1��w<D^oj����S��E�A�`�8�5��z=_�񮣲�.�^u�wW�d�x�M!���R姹��u/
[�/f�DM�A��{V�-�_%k݄��������h7ayL��J����O&�·�v���r !��)��tk������h���a̩=��9g�أ�vX����x�C�3?�~��M؋P�*ߪ�Vp�����k���h% �ݷ�\Cv���{����6�=������1#�M����؋��r^Y���Z%�N��&�v0"h�?;�[����a�B�v�1�O<e��%�e��V��_C�z��f�=����E&c*"D�(�{�{=����p��e�`áW�PU"s&_ �Í��0�����
�Cd�/���ᵰ/0w&d;<?g�*���y�f&%�ﴊ���j�t=_�i�I�|X^�߽:ʩ��R�.�/�3F>6+�z����`Q�� �j�ɲ�e
Ry�E��U�2��J�����wx���l������Ʉ��7L	pa���B����R������	PcI"�43g����/�,
B�&0�ΈՔ�^?[� �y"%Fon�m�!����\?(�`*w���Z�4�)�p'��,�%�y��)ߎ���E1	(��}��g%?�p���U�֫�
���i>�5���%����rrl��L��Ȁ�r�i�Mi������i:�d�R��d�����-�H��I�F����v-�=�L��Z�0�x�?x;w�-��fߪ�!��v�� $%e����h����o%�'�ngu��|���h��ҵ�r��.�ExY����a\��\z�~Z�+�q*��#���{�0����:0@n��c��[E��z���G x݇��^����ƥ|�%�����ߪ�/zg��i"���=6F�w޺xJ��$�H�-��#Y�Пp~"A��`,1G�h�-|@������4H��o���p(�OY�ݏl���k��S��%���l�D�4!U$�����	@n�\L
�ߣ�ʠVDbnĮ@�5�&"��%g�®��`��9�Ku��Є�	�_n0g�Ҙ:�=��,J��W�m	�RIy�H�n�����.�$hc6�v����k�ܳ���
�2�pp�wSo��x�E�أ�Q���~3������h�Sy(N��j�2��lM��:t�F�D>ސ���g /W�ن`���P�a[o�?C �o�8h��;sy�������	9jT�m
g��F
x{4��I��yx:;�������>�~�Fn%�S�[,&����������IWqA�D'�����K��J��3Y�uev]:�N%^
9�W�F�o��+�-6�倘��c��~}�����Vx!r�}�a�