XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����o��Š�]ȑ��6�~i|i�$ˉ�wo������;4�Y�T�=�j���X�wf�L�4q'j��/u&�5��𝵳�T�e�M�ŷ�����q�Rفc��`I'�]{9=��xĄ��p&͌@В���`8��$:�>���Xإ�������k4z�ɫI�����З��g��+<��=ߊ�קyh?��&��[�9����D-��FY�����ʋϗ#�T�TN��&N��]V�.3"�Y�>��{H��[���fGv����4��3�y���U$��J��2|Ǭ�����TQ�CA�اC4`�֌�b�)�W곳i"��F[~�1Ǭ�`�(�ԝ��b����$7^�B|T����G4�kd�Rl�[��SM�]��Nw�g��9�ݧ�ߐ�Ig�~�v�xK�/<�ž���d��(Ix>.� :��ӾE�Ɂ�3��Qz�o�E�SL	@	t�j6#�p|-4��L��+5�~/�46�9tnW�����G�y�7���h>8���y=A]��A`��ҷj���	]��:�7&g��ve�(3�)F_�A��0��:<�'��#��'6��a��JH���'��F4ך�%a�>r��ar�"��zx�Zm;�zR��0��+��+J�R��� �^ɂR&AY	/� ?����7�<�m������o��v��Q��^�r&'�5�<Zl9�4a'-�u$}��ޑ˃��iTn�������ק)���/���)x��VL�@��XlxVHYEB    18fe     880��&4�Fy/|�D��>6�m��iq�'OE�%���o�ƴ�+��(�M��zݞ98�K����y?@�;��Gr�4�,���oF�����*zP�i�n�OU�GڜFH,�����F<�?L�����W��`�>�6�R$��fg����G�7 ��w7��R�;�a�Q��/7` ��,Z�Ju���?�R4	nu��o/|��R�eC,/Ӻ��6�7����d�?웗�4�S %�� �ޅ��\��[��<�&�x�-��u����tJ�]��Uq��n?��!*2�@��Y�a��l���-���F<�`�^:��NG �D{o�����$���D�v&�t��4�C�@���u��UQ>��^��W~��TZ>��
>�!ر�� ru�����|T��8������� ��q���� ��xU��ڌ���v��g���0���ڒ_Y�X���o8ݝ�}%��?��Ә���DJ�&(54RɰŘ��?3����h��\���@�M̏ԓ J�J�I:J>������Ե��_�9�c��'��R鞆&��n��@�e���a톾`����LB�����:�<ڸ�C�<��C@ �E��d9�h�@���4�����6T�@܅
ۨ�f�K"��~.`$����t�n��h�mK$[ˢm[3S�H�&������<���`)��@k�$;���Z�26_HD�����=j66�~j�o6��{n�Mݕ���p�k BmL^�<��J�\](U�ix?��H��z�4�v�S����J���g��S|x�1�~|V>�~�ш�-9��R�2�mFZl�H(	έ���{=�����o� �w��=��-��PU`4�T)MNi�X���cT3�н��g��PD����-@�%���#���܇Z<��3��b��;�Uݗ�7�������)`z�r.z]$e(
 ��\�(����p���d�d�h�s/��!��S	����$<+؆���Z)����H\��2�4t�Y�R5��g����u�)���������S?B+�_��w�}]JG�v?&(��n�������F$�p ��h���hHğ��3d��\��>��I� ���,_9��K�~�I1�K�N����H:��>���-j'I��΁7cj���:��A��1|�zi�Rq7�BG'�PR;�{��y~K�c�T�XLɎ`���Q��X�ה�,�.�3��Z��+�5q[XUо;��KQ��p���J��� �j�4��M�y��=+�//��K�����߮��k��+�k�ͫ`�wc�hy��u~b��HG���1��}swqEf�b������[�S�WQ���n�Vp�Al=y��#�WH�n'<8�%8B�������W���Gv�<��V3<�)�/W�"n��o��TM݀��(_S�*�� �%x�Cr5c�W<=S�e!:�	�x�ɐ���ß<��wz�E�%|��΂[�A
�'E��$�Kf�j�E�� o:�������q����9L�������*ui�i֗Gl����Jͧɶ����Is �Ճd��z�A�eN��m���v��s��"+a U	u���8��?lj�L�O�
'85����\Hq�^���h�L��C�WM�A�j����-���6DځX4�>e�<"��D���Q��6��܍ͭ��w�>��/g�{y@�t9vϚ&�M�z������~��ˠgY��%�!��i���������5Nq ��N�YMR�-�E9AR<��c��XB� O�s}QY"��b�|��r�l�����Aￊ<z�ykWy��T�oC}��=jGs%�(�َz��l(�d�Ⓑ^����Ns߯�]����n>�ߛ�R�̻0���C �Ϳŀa�sAJ,��ib�;�M�~Oo@�����H��q�P_��mB����H�_�|A&��/��s�[&l!�A]��+w����i�]3� ��# ��{Q�&���'�%��b4�P�v�/b��P��,P��Se���ߐ�IwSa�T�̐?����v"�R)��8�nt?"��<����GSN|z		i��z�9���;��k^�HR�Kw�RxHH�Ej�/��ݿʆ�.ȴH�e�qV�SFK�:�O{�@K�'$߄6@