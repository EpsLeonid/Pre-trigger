XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��83b۝�-X��Oe��Y��+���o���jt��eOQ
�դ�̎�G���Q�
,K�xZq�S��@ч�v�q��֨}�:�������c���h\� lj����5����o/�/�{J�Mw8��~��΋����#n�N�}�zy&��%��*�Cܬ�0"����,�MY�Ԝt�{Ԃ�I؇Ǽp/��}h�$o��H�1v�@���� EL�~".�SK�k#�\lv d6�ɗX��%��)��G%��$?���#b��I�K��GS4�g���x��ͩT��%6wqT�Eu�N�����^�a����|����
嫔�%-�+zr��撁v�[�!�o������+���5�X���V�KvQf�5�{���3�P\�X+�A	��6�f���vώ�f�ı��e��<i9q'�S5X*ȃ=[���`J��_V��W�k.6B��y����0r�۵�2�9n�~�3D��S�7�P�0�P���Fb凚���@z}�̔��a�T�!̞�q/��>^��В1��Һ��c���ԇ�a߅y�7p�$Y	�W��ZP�y��ٵi逕�b>'0�����A	�1�%eu����W���l1֋��p|}�M�w�R�VM����~�C�,�)�F��hs�]*ر@P7����,��RJe��5��ۇ? &_a�H؁u@�*f֓��=�l��.�S�
�H�}<�$�0�}���I4Qe�>X�$j]/!4X�R�v�Z��u"�XlxVHYEB    bd1a    1920��:�z��j��֞�P�$G�����3�� ��j�>�`.Xs����&�����L�&���T0�K2�"_���VZ)������+����^<��k,M����LޯE��Z���
{.�?zm1d�g�"!��?28��2�j�q���s����	�:�V��M�>�W���2�}��w��C
�Y�ЌMR�k�5����S�ɍNZ?O*�|����̕�Ę�¶�eq
�ܒ����b�m��	5Xn�e��h��=�d�y#���<�m'�M��K���6Ont-�	��˭�׸�$��s�ec��Y�cXk�?��5�T��p�;�q��W��L��[C}᫏w�缴�	'0�0Fz��ug�d�)��5�12:�Mp�I�Ԛ����o�PҊhCϋ֣v
�H1�����!���+J�{���F�.g�&��-�
�1�Z��XO�C�kᴬT�އ࿪�o��_nV �s~�6�����c \���^�_b�-(�lO���1V�T���h�6�����V폦6uu�,��C#Ez�Y�`j�n�=���W����n=�+C���"F`��nv��Ԍ_N�fI�B�yw����b���.�i��r����3�!~�iF���p���LB��U!�!g*�)GJƚ"�P'+�gq��f�sT�K	�; -Z%�-f��(�<�.6�)5 r3a5BW�TG�
����'8��:�$�#�ȱ{4`3Oz�c���*j��39Ѽ������^*�f��o<(ⓏB����5|�ٻ�S���m�d������_tw���2Ľ'CQ|���l����8zm���r�uk{`O)��`GXj����:�O�+�[��{L�|��/��DX������Xg�f���P��P!4�8d�hB�bht�2�+�!�0j��^��8�01�?	�7���c�ϡ^�&�#M	���I��d8��K�'4-��43���\���D�ە9�ȈB4�=��q�~η��Y��,Y���ʯ���ƹ��H���xrl�bs��u�?���?��C�s]N�/�a9;��3��0��V��0� ߱�uF&[fN3� ��mj	�(��ZD1|��p��ޫ��9�C5��j�,��;��ȁ��f�>�ѝ+r����v��-}ٛ7���F��9 ��*���E���6|ۉ�8Q]H��/Q�v��$W��ζ�9�Q��Y�>���� ʈp����ph5̙���;�9>dĦ"!�=/�;S�e�'3+9���W�����15��W&�EE�S(��~iQ5�C@��� =����
a�k"���$ZW�H��XAph7f�skًVk�]zk��^���@/A�2'�`�7v�̢��ܳ�]��V�_����X��L~�\;V\���O�$�g��*����a���S����5���s�0��40�r���΋���`'/9y<A������K�i�ӥS(��8bMy����0ן�z�x�����s����#�FA�V.�W�����iw�27����-���0�~�8��;�y���K3��̅���}sTM�vQ���h�!�����b�������0F�����AG��,ޕ��Ly|�qQ��(����"�����	��	��H|�X���P��ά��K�<_��F��	_�pT�k�)krt]�e'��c�pw��'�H�n?a�I�����/~T�<E���5?o��v&�6\��T��a�B�=�����I�1�7�X��vp�!�U����UP�<C1A��:�~3OG>��%�ڊ�t"�O�R��ءVK��w�ԋ~��}�'��;���3�OhU^�o#.��S���&bL���|���t:�,"�2 i�YGα���j}ʤ<��>����[��EB�D����tC��*%-[t������ێLl�����@4U���@�v1���R����&�^�a�S���zC	~����e���=B�:Ļ�i��s����g�hn�Zȣ\xe,�'�k0�����Fk�D9wH��Uu��)�X?V1�v��.\��4�,M�<�^��MJ���~�:5n��L���J%�J��S��o�ßH�=�m���֓(����v3���-ZJd2�0��lJR�CM���;��u�iB�0��A����A��C��b�Ы���Џ}9���$��g��P� ܮ�T��wIE�0��$���SB����5���4N\Go�Ϋ;�R;S��/�hf�Ӈ"�3ࣼ��y��!!+���o�F3����-�.����o��B�O�ə�W>�O+w�sL�d�S��٥t`��P` #�4p�h�#<_�ѥ;Y�t�"�`��c����������.3��ʱqJ��ȑ�-xأq��7&j/��g����Y.ɣ\�����U�R��k�0a ��� ׾�������n%g�~"P;�E��_	� ��.ԭ�-c��~�D��]�"���R/�0
'ͭ�&��v��$gN$�W������i�-z�J�����$� ��"\��#��9'�A˜ӣ��O�W�����Jw��L��BV)O��\�I�M�QF]�N�n.�8��w����&4�nD)���|-m�5
Y���'�LmQ5	�f�i�
�+�-�A�/@�<��C��KT}��Jà۵P����J��"�fQ*�_�Y�/w�P(1��ʏ �N�z���lH�?2���~BEvv3���?��c��^η�U��}bջ[�t��A�/F�'�1����=�H��n���p����Fq�Q�$vJ>�lAr��	�e��I�+X��3ŏ@Q��%C����yn�ovpd.�{��3Pϋ���a���q���S�:��5��C����,�<=�Fb.�W9�+C�F��gҌ�Q�Q�^�>:����Տ��_ �#�=��B��'�\�$�S�N �c��c�v&�m�)0(���q���%w�Z"��^�+�6����Ǔ��v#��Zיִ�����-�O�)T��:�t�!ФMs�Y�+�A�vR�PQ�8��}�8ƿH}_ j����
�Ϟ_�o�N2�,4KY/<��CI��D/t*�!/W��")? %w��r��n�������݇��-~}�I�_��k,���'u�-q��9��4�-��) ���
��'z����"�����/��}����V ���tt�y��K.��Ͳ�kӵ��s���h��671������M-n����	c�4�O�g��J��z��9@�� �WM�xMl�u��}�UAN��'��&W�z��&��2b.�k�2�ɛ6���ւ&�7�<�_��?js�W8gtz���|ƗC�d~G�56;I!����F���V�0�����XMI���&kv>鱃a�ŁD1J�)��0Z�blf��!��,I^�[�*���ͭ@��S�lQP4�DD@L��O��V�5p.W�)�����m�:7?E"y��Rv����P��16T�6_�g���{��/�����s�G��i�.�B�e�����'~����[�����%���Sc��j��tɍ������U��ͥ�i6�ƯGv6��Ӓ�\�Y(�I���A(��`�uXnQ� ���(�ț�pV��#l0F?�
N
~�R�~���uF�GN"y�B�����|����&r�Kh��_�Y�� ����d����1�?q����g��m	sz�y�H�"n(�,j��ׯ�+SYe�n�����.h��Vc��-]-��)���Ln|n��:߭B�B�r\���,U�L��e?��b��QĄ�JCs���*?��=m4��s�����dߨ���1�%����}�G:�O��kf������\���v��!���Ú��Dn���	�GI������G1l[��As -�	$=�N���-��e`&�4&�.K5�5 f�����9����;}j<��1��ӽ"p����Z>y��$t����H�q\CX�2�G�f?��Zf�WdH�ڶ�W�p*cX��2W�j��@Q�i_ߺV��v����nb�v������,s����CJ7!�2K��f����["���nY���[�����_Dل985!ޛN�?uӽ�_g����J�Í?���`��sf�x�ޱ�wGבE���/�mbA2�aX&��>��,�rV8��'#0^�?�����}[�TF�{��O���LԢNn�� �\�^���ˮ*�u���Vr�L�mEFץ\b�:�����f�>�̄P�Ř�����h�b�K�"�������� u1c��^���U�5���^Y(�^��v>&Dk���ϳW|X^t��o2��|��(
#%�]�}9�{8��u28�i	�yK*��\Q��K�)��y]�"�GGT��WN���Si��"�A��:@���[u��!�ҍ����`	}!r�KX�#u!cb����/�%A�_��5B��N�S�ƿ �̮���ݻ��]{��0e�^t�Y�y@s����	j�6��`��@���~x��A%�9zC�ӷ��$|؜��7&��=<�&JF/�"H�#������/z��d��+�P%)�f��dFL'C�u�f����n�w�0J��7��z����ޢEu�Q&�B�m�5�j��ܱ�.�����D���D�2+C@�#v]kR3���%�"��Ye���V+��v��O�Π|й�X�	k06t>��ʩ]�^�w<��'�'b��+��ye�x�[wT�}��q`��AT�w�p�3D�z�/���&����VH�)1��|��{�1!W#�{�����pk�Vⷂ`�E��9��	�|����<�C5��]b�>�s�.���চ����C���}7��dӃ��s��
��y&�.h�E�3-M�n����j���)\@�o�&;��DD|��`�gA;�Z\9�L �,���J�{%��ao����X�w�DN��æcf��xi[�R�4�>dq]���@��!�ŝK��ău�Cmp� ���4��|,���������9$..q�bq��G�\%�҃vQ�
]��gd��Ύ<5R����̒Y���80�/�_��x��ZK���d�8x+�ݛ��W���n��I��'*�ybFT}!���-���~nf���Y�˹��ŰJHf�Zu�x�U�^��e�o?P�<�8Y �}��@T.��q1O@`U�� ��0֞AI��b�v���:ʺh�=��A�K�##�wH#�,�Ǳf�R�M��,�N����D��%0șb��();7�T�?�/���N�f���7�=�����*Ŷr���F�������n�3^ Ȍ v!���0����pK͟���S$hTG"+(!s_4�t��hHn����q���r_	�06o`��
��*a|�N?:4�p;�BH�\Ӥ�B'�?�)�Ir��	R�V�Oy�Q̽u���67,�uӟ�Ɵ+&?�Õc��'m�D�A�jh/�]9�ѓH����~Y��*��v��#�dF�"�3ZD��؀4����ٛ��+m�R�?�k2)}N��'�� ±����H,��}�M)��
v��UJa,�lT��r���_W��@���$ @��Nxg�jb��4�2d�K��,l�H�=%4i���K���j�zn��.k�CЗ���}�Jj���*{���ѿ|�~_5��~{���69S ��/�2������xST�B���>����ȃ��-'�=�x �;.K��	�Y!��b�ܔO��I|�葶@���[���C��cP����4�I���򯻨�p�(���V��M��B��#�^[ۣ����^�I��.Xr���ނ�<og`�G�1z�l�V��?�����V���SwI6%�9��e?�NJ��ϡ���~9l��^?7�4}��r��K��|����$kIE������jm�����?Ó�x �Jjqyn�ʕ}��j]&��&Q8��]}�@28�3h��)o�`��<��֮�,㣖��2��;Dn�9��N��_��M5!UNl�t��I�Bʧ�$lH�0�e��2垣�A�Q>/���5�p��j
�M��)	o��t:CƝT����ټ>��Pw3U�zL��!���	��ZY��])T�:����@�E�G��=��kىcf	M]Bͺa���s�fJz��/1i�?6Z��z��#T>�l!���;�r��\:�:+�Ɛ� 5Z�$��>��ڪ�vr�Б¹-�� |��4P[8���}����
;�1�j�u��E��UZl$9?�����F�\#��%����ߓ���b�=ȻA5Q��S�lr��1��}=����a)���M��l��ts������KnwJ綬a�1��56x�g�q