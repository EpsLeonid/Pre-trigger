XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����
:��m�8{�p&r>��I�W�;�1J��XW�T*7QC�{x�R9c�)~Ȩ*0��+�)m�i�7��]\�J�8��[�U����^�OIŅ�V
R�%����90��&oR��g��oޗ\rzP�	�ODӢ6�av��������x1��O�ֳ�<��\t�C[a!�H{#�РCk�0;a�m���4��/�<rU��|6��x�p7CC�Ǽ�A�P#Q�OĵcnexDy��J�2"�:6-mp:0��d��� ����B�\Q�X��$��г&ԧz.eE0��s�"d�yn�M&VT�&xF�L�"��v�RH�����������B 9�'~95�D���W�z(Ĥؖ:��;~9>�cq~������L���W�H�#R�%SL����B2���/��KA@ѓ������yF��}���o���6��Ʋ."��q#��$�ɇ�ٺ�D7}��
��Ug�@��T@q�FI�A�(�b,�[_���=��b������zǙӌu\�z#;ü㈇�M�`.�V��b!@��*k���4�`\`Y�ʯ�M�Cʉ��$
5��8�dVL�>�'���C�i��FRh�ؕ}��D��T�T��\<&�]10�"L����� �{�0�Dt�1*_�Ƀ�:�{V�Q���e��>g�	���*9f}��P�=��`6��x����{�i��<�@X��.��M;��I�D��Aߦ@�XHm':L1:�So+��OM"G�B�r��N%GO��EDRR�ʊƳ��a��nG���@U���iXlxVHYEB    bd1a    1920~�k�k9�l�D����l*� �Nl���'�m��>�����XM^�eq���0���ztfEeىcX� ��|�gN]�����4Դ�W�ck�x��8�ꠣ�'�)4�& b���F��d���R�N�����%-:����J�Js����N�G�~C1)E��U�>_,'��"`�7眝a��Ӳ��R�@s�,S�l����7Rw���A��P����y���a唠o=J�3�+/奡V4����^����2܆�Ϋ���0��RA�8�t�S�V��d���}�ƍm:�,;p�gbӖkj���ST�m:~RK]�g^��C�td�}+����?���,��X�\C�1������V�K[���&*'�Dښ���Γ!���V��lS�K�ګ�SN�h����[@�߭���'�4$$�r<�m��v�KQ3��1㸝�^n!��-�'��"�P��"��<:2��r�����pZ��o���G2�����V)�O�@z�܊���vѽϡ�W�T�0����������S$��!���+��?�<�u�;l�Ю�|�Z��}���-2���� UE�������K����9�ߺAtb�޸'�����ZZ�peg����%SV�Y�-�$�{
������O�	��58�8��=�:r��M��+�0�M���g�rq��/�����0n����YK��F=fN�38<�v�����H.��̪����w \f� ���Y��I8�W?�)���w��e��>r�t�D�����&���(?7��H��_��U]�!z�� ��G&�� ���+�i��$��b����{ku�ZtQ������ݥ��/��&��J��6u��L�N�񏌞�&�с��?x�$q�t".�4� ��k��[��9ѯ��:�u��I q���bu��	(��x��OU�pz��52�7��&�3�(�?���%U#`��M%�_�ü&�W�Hs�6㚛"��;:���ɦӀ��X���!�r���ꐷ��>R�mU6�]��{�W�ӝ~ �<��Ƙ�-�(���C��/�w��T���㡠�J�.�%�H^ւ�_��9��^s`,������h�v8�V��������19G ����#Ǉ���&(@a���=��K�WrB�b1o!Â>��M,1�˕�F���.+���qA��rY���B�7s,��$���vᮇQ�k��췘��]JgW���*@O�+Q����f���Ow�����3�hsP�{jokNf�!	��9�Di��F�
ё	��Y/�"��F�֌���/�H=��\Z���d��
��"����g�� �P#:��|��y��I5BÀ��C�����<u��-@�����Aw
��g���z@G0>~@yǒOC�yH�dG~Ǚl���J��ji�?~���X�'�p���(訧�$��(�����EO8�+�h}q��/J��mT&�%�˥Z}���ɬ������JOE�����k%�ڙs��l� C��c���	l���s���ʺ=}�e���U���NDZ�Ā�P�3�ڛ���RDՊ�\���@�Z��B~����K�⚽�F�o�)"~�15fZE��P���Ix�\�e�۔�3��(Aes��F���0�Bظ�ْ�nT\x��t�eV��q<�3ȷ:	��8��ę4c�PMr ����o'1�N�`Fhz��M�U,�8��mV�� �8A[������/���/�c��^��?O_!���.����ݚ��+��^��E��G��Y��ب[Ɯ]�t"�2�7�[�N�a�7�"EȪ(Ffώ��Y���2�_r��u����G���?�L�OY��C�p4?��s%�S
&v-[��T�����'%��C��>T�s�-D���3����/ {��8�a��q�e��t��,�L�����؂�XU�hت�*U?p45�I�@�v�O�T��/��[EAk���UҮsȺV�B�;>��¼���N硥nܷ��E����B��i���)�G1���^m��N̋��OާԒh�V�x�X�%R��ÙQ?��K'V�݁�G��/��������Y,��V���ߙ����;�xw<x-n��Tt?_{�8�͡)��!��g�p~V�=[M��C�/�Ψ�Q�~$*:�R{ݔ;�%��	�+��Eέ.~+�O��a����l����$�g�p3W�5�����*�����
����Mqvd��&�u���a2����/��m�,5�~б�sa;�����_W��z�,n0�.S���f�x�|NѽXL^Iι�c�(����α�w8�B��	�@]D��"d��C�u����%-�{��Q`~����]K��C�Mb���pNKy��TK&T�sm�NP�ĥݿf͢�?]���ou��0$�BN�i �T�/n���3^LH�%�rm������[�j�8ɋ�Y��y�>�V��J�2��D�Z��I]��6�����P!�R��9*��{#ժ0����3�։ X� �R�i(� �z���	dPy�^=��}��c2��M������T�>[������ť�kH���zZXh, �$��f�qg��x�hJkD$�m�~��Dt�$[L��1�|&�91������������h	���d� �C�+���E6~,P#���Sg�>�o������(`-
Vk��H�r�l�P`��8��6ɢ>�ϯ�[��!�{�?PݽY�L$�:	�U���~�E}&�U9J���(�L��G����)*��+f�~Wm�w�uE[uCB���n�>|A�WgW$���Hz�B��@̴�,Oz�B���"Mʶ%1�&����_ol�j�v�NX��`����F��niѲ�`�CKX�/Ƿ;Wx��s��Fmo~:U>��J �r�+��_��=k�^1��oiY�����q��\H7�z��)�g	���$Q�9a��~<�^�ܣArp�a^<N۶d��f1��h6��~^�ѯ�?�C���T��.���2pw�ó���¸0dm|y��"�x�ꊕ3Y� �MoAU�Xk�G��U[9"��=t���ZU1�n;No�О˰3K�RRV�ΝWf:���ƙ ��Z\�^�]�;@6�f08m�=P��;��Ӗ�T���+�k���c��s�u������u��u�]�e��V�1[�+0�-Қ��>��K��~�q�m�8�����s='FT	���EU�@��n�?��gW��8ޠȹwA��4Rܧ���)Z���y�����l�;�A1�������w�A����@`x(>�& 겴r�ϔ/]
�u����v�v�|,&��:j�dG��R��g��yl5cA�&�,翈a��kY��{%�5���	��b�O��� v��h������
&�G��PBwK�m�Q6D-��:���Io�q�xT.��Ogn%*Y�#cʎ"m�uho� t]SN��HZd�F���:qiYṣn�Gi���n�4�2�H�%�/����e���V�-�g�����{P�@�<܁5���j<������Tg�M�D�.�����\�S��\�!_f���x�L}�|U��,~�U���V��_��%=y�^��
�}x�B��IW����l���T��m�rV���<l�S�P�w؈��Ž�T�v��F� �U��ppɶ��$�I!V�j�9�B^�\y��K9�^�#�����!9ބ�����������X�֧��,a���"0l��9�]F����K�.�B�j�<�U�G�j|�M�n##|�FV���eV��>7]H;%bO��2��O%�t]��ݰ�do�9_�v�H_)/Ru\����,mk��Lm����l掵��꛱Y�o���sT�>��:��a5�
�(Kwpj�.�;t�����9����*M�NXz�<�U'�W����"�:�5���Cϙ�\����B����VѨ	�ciL�� ʗOci���S�_T^�ƫpq���4���MF�N;�Nάw)�}�U9I�X o�n���ݙh��S$�;r*�v!��@{�S�\	����4��Yv!�I+fQ%b��)�[}&�$��䶍��,{�#�U �p�,-l<�Ĩ����^�$
g�D�&���*�������6} �<&٥�w����D�x�ի��ȓ���]�� ��B/� m|{[�5@w�x�Rf��[`��80'��L��'�Z���R��D^��H�P�.�V�u����\�J����*��^R�� �渺����M��)HJj=;H�ι>ۉ�/M��`Y<��=�OXQ�T_���n&
{���,�Lڃ#^뭦WJ�Q�?�z���|�rZ�1����x���D�[�EU�|�K��=��gR|�- �a�tZ���B�?C{��[�>�H�q�#�|������F�+�<]��b��7���P�8��>��/�{���`7�߲��aJm鮋6�C#g�D���āQ�F��7��zъ��W���:<q,�T�f|3Xp7 ޅ?kT �*�xݨUgcG��ŀ[Qq��_Gr.�=��h RGO	n=�9�WA�}]P���7�T!/�krp���W�O�g��X�m����\���]S�̜(P�)��Nv��9SpO�����ٻ�~�`:��^k+�輺
��bL%$2��W!o���,�O��a�Ɋ�������aG'c�߂�$�?ٌ0����_���2�,h�&�����;�*����� [�ǖ�iZba �yD�m�5Luި���>ʶX�h,�R̃+7{�'�]�Sb��a{Q�AM�2�:y(���D���D�#&�M��m�Ek�0J��tyɹ�ށ}��3�����D=��5�5�e�&j7X��`�x�V�,�nUYC0������[���8.�SJ)�m��k�d��B��\d�;�6�Ϩ�FqQ�G;[<���9:����i�y�T�7��s���v/7(IQ-�)��[��wa1�)s��欐$,'7�8�He| !�T	H7Aا-!8r�-(�ݒ��X+X'��dn';*!�w��",�`�.�(N��=@�cbf���$����uEݤs-4�LAu��g���~���ƾ��gY�g��9�K.4��Q5��8��mצH�F��kK��*�Ω3����Y��R���-G�v
��Q#����
�)��ܙKm���ۍ��-/�6�}nm������S�~)��DhN�ӑQ��_�a6�LC֜],��Z�"`�,�r�gY��+���V�Ie�8��*([�&�$�:>#��>�������iQ6��c"彻vݘ�O��d\`�=�M���R�0��Pw���墴�^�r�~�{�p�T��,M@��!���$:s��7w���ı���w���zB���������K�o�k�9����21�XT�TS|�b'wk�W�u�R�����w���FZ�K�o�/�i���2*R�k�4c-	% �^�����K<J%��ȫ��.�8�! �Xȥⷨ��+��sG�(��ە��7�G���b �Ye�侇q�?:4��ĥ��܁�ĤB�S���Z2��fc^ޗ.b��u$\H�v�2Uό(�j�Cn�Ww�2@��ڔ��?�d��`��� �XU�=���RF�>�X�}��/�0f�~x�@�<Y�!�p��؛M�0+���(`w�EӚIO��C�_�qݫLD�kf��o9���w�xe��	���
Ua,���dU��=��fS��fޯ<1��(��7���/:��6M��'��2�DG��y�J�g�Yzm�Eќ}W�D��9Q�T��f��Wy�D��;�\4���}�-���?s��9��H"�m7]sf�Vk_U�i,F�f�Ah����q<^��8.0c9��
/Wy�W���0�I��;�c���+��6{�>8��aV��I��_خ�#6�Z���L�Jj����V��z>�N�
W$:���C�S8v��u�ue;�?X�,4���h��\�F1'(��g-�T�]�.x����:�pw3��N�E=��0Ճ���cCϸ�]"[�0Y*�U�\/_�Rz�'������Z0��C�V�)#�i.���%j��Z� ��e�36�D�6dB�Ů��s[?�kp�'�8��k�(r����x�W+@8��N���iV|���j�0��\� P�j�k�u�0�Ќ������Q+H�df/cQ�"Tk��W��T�}��k��[KΑ�� �p�^��^.ec�$��'��&i�*F~E���WW���z�1�C�#^l��0��}��9��L���곛b�ɒX�[cB���g�]���w���"�2�