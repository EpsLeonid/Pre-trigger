XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
���ݧ��`uq��;9i7���3�C�]T��J���DίE�,!P=�"$��/����p2��K�ߙP���v���o�m7��~"#�l�8�r�:�'m�ǅ� ���`
�xW ~`� i�D|�:9}y�XE� 'CM���؂P�(�#o/�'7�2;.����Ʌ�XA3{6v'��) �p�Q��᷉���N��f���5Zm!��7����m@Z/�����*��[�9�V;��*JQ�Z��t'�wk�ǂ�O??��OhQ����0���eţИ)t1��'�����U���'��7��,ì�k[���\2W:���7ϩt]�k.,ί������^���̜�A���Cg��Q��� 褿��8�7lZ �?�OG�%��}�l�㛎�hQA�:�a��t�I����h�z������-��;��R�ї"�^�`]c>uk09um~y#���
���ؿLA��W�v�W7꬚b5��w���;���~Ƹ��௒�&�rciØjm�������6�����+�>�>Ȅm�x ��Ň���7������=O�iB�e��� �K����!2*W���P�q~�	����†(h_�x�y7~�ߞ%ޯ�h$��fgp}.��,�?�Q�`��X�VRg)S1@_}؟Ts5�^&�
V<q��Cn�ǔ�>�=�u�����F<ҽJ�]���E~��U9��P�O�(�Yu���C5��E�и7T�h��D�\:XlxVHYEB    2fbd     d20���>�Oy_�����.]^�,oیw�:�Ѷ�F�3� �5����vϒ�5�'ܤȜ�̛�|2s����1�Í���W�����E���7?������]�)矝VS9��a�oR\�?>J��L{�b���Ư�J�.��@^��(+g}s����}����}�7�dP�F�؇�J��y~5�����H�4T��ʛ3�d���whH6!h�(զZ}�h��~�9�Q�7����w~3�<?f�ܔu���`v�1����V썫��
n�Gyŋ���������m��w�:�:�N���A�cĿ�[�������@�@�q">�9xC�]3̻)n�C���@r���7������E��ހ�ĩ�$
�A���U�N7�\�z��'�0��v	��lݝ��N��(��T�D�k�t�H"4�R���CQ�쵏�w;Y�J0[�|���#��[���cl�m�2xL����1 䉱8/ c�+c�Vq^߅�5�jTx�̝P�%��#�cE�-�[N�zu��pz$2�[���ֆ-�}Bī�����+�eME=��Mh���:z��VAC�JC�4s�԰�B��q�>�ym�n��Q���Z����� �_{�f� c�$D�k��E�I�M���� S�&(n[8y�@ ��g��ؤA�~0���qJ�Ud�MVͿM"Khm��*�hH�V�@�Ƃ芺m{���H�����r�W�ӎz��L�� ��X������_L1!�����
�DD x�`��F��/��rҝ����5~[�w/B�V�#����'�>wu�)){�0�|ût�S�O��-a�z�����[׿�.o]���X�U�OzQ���#Y1���O�^k�Ϡ���&*t�EEI}W]F��K��)up'��WKC%���&ŮO�ovGa��L㰃�'�c����N�	���(Ս��2�[�'����6�{��θ%�Z�o��\�?���ts�nWLd]��[=���`�z�Q`@�ť����-�\�PV�����|���u\�R�'�ָJ����\S�E��j�ԆO�#��"�F� E;@-j��q0��'X���;��܇�\}�Eg�@0L�����k
)�.�*'��������Z���)k�R������4��9AQ�n��z&&��w2�%��ʏ��͙SF���%���4%uڢ0�,��ݨ!��2�2L�5/Q	�	?mڦ'��NI�6Ζ(g]�����Q�������*��TN�0��=q�G��[
I8��K�&�����݇D4~�����[���|�}��߷�/�:"����2����O�����0�ɗ@o� b@H84}�@�ASZ	Gݤ22�	�!�W�¶���UY�N�g�u�W�	�B*~�V�-"�P�+9�Y���dj	�Ou�b>����a,�tQu��#o8��w�1��@����bG�XU\kd^X.�`G{�.H���@�t	h��	ZD!7��xf
e�w�T>c��Y�	��f��@��;�XW��4��{�5@��\T�ǁB�v�̾X����0���~P�V_��Q�%5]��e��U/��_\'M�s���Hb��4C�몡x)�anr��l�=���ەv�+��V��pBQ��C2_uQ�UnH���.�Y?{�LP�����A�g6瘆L:0́ҤFq5�Ŀ�+uγ3��.*<m����P;�z,2_`���V����� .sH>ε���Q���lN�Nm.��d�C��I��| �h����~u��W�{��B$�ԡ�/ڑ��,�5z��g��e����$->w�KԤ-�0��G1��zؙ�� ��]�n��q@�Qu>�%�А݅�eQ�HvH�Q����	䆬�|䈩�O0�X�3����o�I5{���rn��iu?��#�\
bA>Сi����e�W�$�8�T�+_��%\f����)8Ų�.@?���l$1'!��x�,�4w��/Y�ثzt���<���/�S?
)�f��oUA/D#�����2���O�`0�6:9-x�P�{i�X��ZҺ��,�Fe(��F��A���˷� ƃ�/�������5�C\���歠1@Z1:���۷j������:��q�W�6���7�JW�8PD����*a������*<z��E�y��Y�^����ɳ��V�O�J.u�n=�A$�6��5i^�@�WEG�-r3����z��_&�+u����둹��̼����9��^T�e�b�YO����i9u��C{�y�/阩#�����5W��2�����j��Q��� ��F(O�-P����t���&�:%BQ��*�	�)�1��c|.��LZBS��P�i�_�W���4�z�
	=�GR6�.	݅�β�Nh��pf�j��rU{m�2�CKU��W��;h��;�e�2�,WO�$�{�i��A���Ln)��Z���o���fy���81��;�}t6Hɑ��}G����t#1v|O��.I�qEF�i�zcy�n[y��u�3j���[}a?%���?�"3��P�l�8�6�n���_Η�)`���_cZ�6�S���&�����e��ɣ�-k�*����C�)������@(���A�2p�|��L��!@BM��z/�g�J��#� E��e��7����;1ڞ_c���s0,�*���_������9x=hB�X�Y{\Xf����H_�B�X�\��vL��ǧ'�mgDB��� A��a)v�c�s����yK����,5H����C�����7E��"�3�+��lZ%����wՆEj�ڛ�.��'����l��a��.$b�T��o)V�m��7���y�
���?&��}Ȱ�?c��XB�4y��lwϕa:!��偺����3�/�J�:��t�"Jg��Sg��F��*_[o`&Oy0����Z`4و`�M+YȤ��;����@UCo �uP�D�ԩ� ����}�S��qfI��Hf��\69&��f����e*H�����@� N���OdJ��`�e���ǫ��?t%�c���嵀g��m]�1zSuB���^����IO�*�(�:_�T�Z�`㶺de��	f}ή�V�hf�M#Rz�k},Jx:���RjN���2�1�"Հ���͉�	��4�nk�М�a]֡��v��a�|�j�#��Y�e�[��!�D#�CS���c���t4�J@LWi)��M�'B�e�R��\ͩ���m�qt�SulPj����mA��	[5�����'*����Wְ�h�:�/ʏKExnt��+X@P���i��{px� ���)�)��_O��;�J���Z