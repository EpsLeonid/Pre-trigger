XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?�=W�8��­��+� UN_מ1�|��z$��4O33h�6���#��a��lދH.
�������b��|Kn�G�r�8��Εz�D��e���)�	1�/�Ә����m����u�c�~�����k�U�6��&8�Hx�`㎿�&�\hL��M�B�A ���%���%�ˌ����'�X��^�-"D� �Q��>�<gm����6��m��������q��e�Zq ���^�#�&����P�t�2;�)�\��%	_���TGtvBZ���:3����Y>I�~����V�G�i��u�u�t�&� q�	_|Y����f>7 ���嬓��R�۹/z=O�[��IT[cy����r���VÈ"{��A��\���w�])�|*�O�Qˏ��QPD�>}Ԩ�.��./�����2��{�R,��"��Ce�z!��j�2E����ĉ"����LiڎW5�ɤ��<�$�J}E=R���0V��K:���~uh��fn���^锿�G��w�� �d�D:��x���.�	'"����d}^��p}���X��*�k�\�n����68ʫ���:8 �=������~�M���xc��jn�0�d��p���6�#�,l�B;�. @"�9~x0|�����m]������]�;!����x_��\4H���a4�ܗa���v�4̡���k3�/[}���GhN��q���V$gO�x�����T;TrOY��#j�c�tA�������?�9:��I�XlxVHYEB    fa00    2c50�ёDa��_�����؊\�.Y!��d��*��3��p��-�/"`�7Z�־�&�-	[eE��Q[`%�BL�e^n��}i��F1�uv����&�I`jH����|����E�Y$tY�Eҕ���`<߾�Ӊ���˲ӳ�������(�c�F��=r��#��N6���o����<~�R'�Ո��Ĕ"A�!�C�c!����,�	ATj�������6�H����2��l�	�]F�0�>� �N��-R ���-��`�CF�`�g�mʛ�H���>B��4�\W ��[lm��͕�U&V-����S(�X�pL~mo.<u�f�]������q=O�<�N�ʶ�S�n�=��u�U �~{�|#�/x�U��<��ۧC�]-?�٪�Rx|K�$�,��-O� ���Ӊ���煎�����eC�I�Ցo_$��� 	�
�6��T�	fU�O=5���8ؘ5��*{h�D�*�!�]�#�r���Ů&���[�;������`���z��LJ��+��n�k?�.I%������-^:�/�N���L��;>�́fΪ}((��5�E�X%8ru9@"�j�0�>ǖ�4�f����ܦY�%�� ���[z1����������:�UA�}\��@,�-��9_:S~䐵�Y��;Sx���s�����Q��n��|�@[ %�~�_b���2�aѪ�1�>֧�*! �xD��t'�C�樚�$B�� e��9$�Ɲ���4�u��F�v���������hA�y�O���r�:��d6�b�[��hb �-��+�T�"�S[��$)�͔�ߝ���	,�Ch3�B�?��'�`�t�E�@fh<��d�ZB7��_���O�')ɪYj���@Q	�{r�ۇa6�J�t��
��n�Ư�&�V#��3yVwQ�M��Ja�U���1�(Mi4%�W���z=L��o���,�L�i����ޡ9�i����A��i���.���l(G�߂~
���N��э�~k?`��x�t�B6�|i��>U/���@����-����^�������Pl�`����2Aa##�a��g� ?��<�`���5n��+�R�~� ���v�����w����b@�u���y�Kճ�)cʌ� �t��\����K^�$_�@Q���`�̮ ��?��>:'��P*�%Z����1��#���F�o��OY�\a�-�z�﵌{Oע���B	�\@&"�y�R4"�=Te_��!Җ�
���T�Y��_dc�� ��l�rB޵�rpa��{���@������,����ӕfʲl�Ķ�h��0y7u��?Q ��=a?ރ��"E���^?�~l"�q��F5��_^\�}7oc8/d�R��ܱ����o��]�c����w���g�&���}�GAnŬ�'��{O�]r�ˎ;��Ux�%�#�q`J^.��~�R�$�
L_4{���f���~/-�{��*����t"bR�����D r���4����'��;��	^��E�Q�>�n�G���#��![��h���,q~Q<�MƟ��&�\��n��]��qp���]9\l�7 �a���Lf�*7cV��F���F'ѩ
U�$A�;�T��H�I���)�Xר�����߰�;Qp�{՘�ሎ��vܷ��KD��w8Wn&�U_u�SHp���Ḝ���*����~�R�"\��Z6KfZ��a�ETB�����|��V=�*�����%ykv�����!p�U�A�B�J7RB�F�E�J�6c�����Ʊhbț*�����7�X��T=i��'ű�^{>N)������1%�a��l�$3b�s�L�³��#�i��u��"|7��0D��p뜙���Yd�تMBC2��>*"N�W��}~�C�`\|�
��u����m:����t���O�V�eE/ �8d��f�P�������.��7�u.7�1�Ԋc�>}�.c���M H$�/؊>��A�;��k2m%����ئ�zu;�J(�o��/>K�]}����KΙ��и���e�^J�=��ի���H���w�I�o�K�B�VV�M��h4�)!���PK�,�I��M����.�.��1�{�#(�{ي�9=�&7/[^ O(���/P]m~؃][��:/d���� :��{������5��8.�4"N\�N�c��>��9�]sk
�]_�u����#��M����蠺���/tEȢ .��d�r6�Y��h
�2��U�F"J턟E/ŷ��M��D��LD��xi�T]�ުt`g
}^pa7NO��v���}��A�A�;��� k�0%oki�B����m����SӁ支��2m�Cҽs>f�h�������/�U���2��O�>�Ӭ.�P�9?xlG��_��]�5�*��k�^S�}�C�� C�Q�8������ZJKׂt���.��Y���Y��g ���R^�u�8H�ik����t���x�O;�Ŏ$�R"=�u��A�	(����J��>�����T����+����1N��x�H�-�/�DP�s�S
6� %n�
Hr��J�K��)3��9ܺ%��̆H�i����{�o�&���C�Q����h������f���y�.ڌ���p�#�!��C� 0�8^�,���.��"P��T]��\�\q�E�P��4��.D=�u�+���v�%npp����1�RAyߖx�V���F��fF��7UX�%~?�-��1�)�{6��(���1|{֔�E�xL�9���q�oQ�8S�;�m�ȇj���jPР�Yw�}(���r��s#	��߷|q�rQ���ڇD�³)�m��!��L�z�X��S:ogS^9�����0$ݳ[��Ԫ�e0�-��l�F<�s0~���|�*'UPAG)�{EtD���Οݮ�o�j�
�ù퍿r��L���L]���X*"?��H%�����B;�i�G�?�4 �����cT�Z ����3�B����~{�xx���,����L�j0�g��{�,{݉���hg}�[��J�X����%
4.�
� Ƿ�R|�N��Ì���K�ҝ���|)��WCY�����ġ^C��c� Ϝj�XH��Ɛ+�	zT�UUh?1P1o���+@�L�����X�fn	�Fr��,��$��AߏZ������v�Cor '��tc��yiO�5�Y�������ks.��>��SL���y[u,����9j��E	�d5�K�YwV��9�a�6�e�(�Q�x�����x��)�r��_���!�a��fʙӠ|�&t!�k$q<�K�W�&�Xt3���H_���9���o�B"M~�N������rY.���ȸ�\�6/��"V�U�u�͡��^�S�=�������j�ܬ�M�a���W���-/����\�sA�* =�Wd���u�=64k�NkT��*]]�����.�IQ��色\����tg��[U!��:g�})t�4��/��`�8�'���w�OS�wA���[O���f�D�	E���*v��+��燰���I�ѝ��Z�J�"�U��@�e��,l���u,b�v܌z��qt>�B9�J��AM��hXߧWxX���5�Z�n�(3�^�c0W3�@�����d������[�_?�$�M�Ε�u�	�7�u��F�a�u��[�:+ ���m)|�m��Q�N�b�A�f�*S�>
^��z�(�� V��1g�Y%q?�	�ce�!L�fc�k���鐎��$���?���H�����,�CD0����&�y	��!?=���w.��+`h4
�\#_��M��G��M�eewj��U��~���C�/6ԕa�Fd����!��v���P|�< cv��Ho�@|��h�:�X�><;�W7($r��l�v��)���Uw����J���Y�*���7I9�B�'�azA����V��K�U!�v�
��V�1;�i[�O���j�t��.�WCP'�T<��[��l{g�(���B��6n��B[J��gj��Դ�l��� ,֯9`k���֡�M5f�8��i�X�T�Q}�O+���?���U����G|
�eD�tea��k�8�t%�f�8\p����f1vw=��l��۞$�O���S����!�ؾHCC��(t���F���AT�@��g�Z1�g �xp�8Nˍ�E��63��d0��{�S.�ՑQѬƷ��!y0�Y%�Q��[A����"r�blU~�;�Y�N�fw-�HI��(���6W�`��c�YB{��\O�c����{Q����y��b�]�|����V�}f,>��=�tZ@���l�$(���_:��!��q��ְMdD�ٖ�@%�اu��k)��G�ͫ!E␱o���������M�ǰ�9�����M(��a��ǿ�������^6�5���B�g�!"|[�e�xr�-�f~Q`��o�5ov���\X}��$��ں��}� s4h��D�ǖ��{I���6*���:�`���~=��4��{����P���~�^�	0�#���E,z'E�HE��GKU�R(1�z�&��䯼]r�ۛ'�pWY�i���:��+t������j��a%�ך���T��	�W)_o�a���E��^{F��W(�-&���oN����@p~��%��[��Չ3s��&?L�~�|76��`����V.���]*�l�U^�>��u�r��=,�o�~�ZB��pp��X;����y�5�����Dr0n}/$h��W
K�% �xf}u��.MQQ͋�K��������X�~��j0��G����k�����t�/-��9j���Dr���йzqЎ[�r�������#�ߖ��F��d�O����I��ߦ��$�k�s� 0<:E�T:����8����.F;$��VB���:�Z��;�'7+d}�&��L�{���v~ѠM��e.��TϤ� �Μj���&dP�јi�f���ݸ�q#bIA����W�|)�F�$�����0l^���WS�R�����fV")]錤�h�j���N.�~D�܍���{G��^��C�i�g�~�bL��(Uq,aΥ��ȣ��;v��z`�>g�a��S
���-	���5/���`?:��^��T�<{���8�Kl�(U�K������$������qf�ۛ���T[6�a>�`5s���3G��k��a6Q��7"*����][�9�&��S�Zdn�\���x�K'ϗ5�S���n%��L\��"�@�*�!0��b���|���@���z��*�������BK��z����=�W��<��X�y�8t����\�ȏ:��]�.q$n��5�#�Uv$��FR;��.v�?1!���u�T�JF�����ꞙ��4���<V��{|�,e��+��w��,vA�hpX_ G�緘Ovj������ʧ96{�LO=]**��K�\� 1��u�D�^,������H�B�,tRc�;i�w	Ny��,*��r�ܤ��'`��Q8�:�,�2>IL/�4�z���ͶG��PR�3n5؆���F�����p=���2��oK�q���ԕ�����}t���~�m}�0�bk� uL�u�h�g6nZ�_�0U�Hu1U�IY^�"� �8�����qp�Y˒0��d��x=|y�#����M�	�H�5/��2n�D��a��9��E-�C�����~ĥ��qx^�=W���F�Uw��n|v�(�g}T�;��W��K��p���p~*T�#'���>e�tl �(d肫 n�#Q��HNe2"VD��Y���J�[��)�������h��޲��b�-@w�6�0X��y��E�vw1��(k��eu�7N�zZ�u���?`���� `�՚� �#�D%�������y�<�&04lfq�Kx�"�A)<^�O�N%��\�yL#���Δ���A���Z�NԂ�i����$t;����mo�w���0����b	�pl�'�Ôj:=~\l��Xw�x�ŧ�!�`\�(���&cY��W,����I�r�v��U'dʧ��ɩ�#z�4�?�q�'�G�w.1[M�p���b��%Le�V�q��A�6C'��_1�hшl?�=xRڼ���+�ebӘ^mH��#��]jX�z���V,
�B�?1.ɣ��aȎ^��#^�E#�P��P��ڑ���Ձ��r@a�36lX����;k���ܜ�J��z��br�n��?�5�Qm�	��OE7X�6��3����Q�ӳ��:§_�4E,�Y4��Z���Z�=2[�w���C|�h�N�� v�,C�ϣ���S�`r��+}�:���q�nԖ�z`� �{_�5����?ד^�ChGh%��"u��� ����r�v��O�j#��u�!
��0���L��#�i�c8a"����/�Ԃ�,��u-f΂<;���"KA��刀�tM
�eX�%�`<���1�Ó���p�|��FAUC �vm�� ���A6�S������?G�ID ����.6^Vw�e3�'�r�>���2˲�1������uzTNy��J�ܿQyt����#:�+�a��F�UV^n�0�^'�������t����>�Aضy�t��O0�Y��E}m]��=��M@���lVx�P�`� x7��_&B��Dsb�%����D���o�6�MN�:t���x��%�'$��,5��wo�H0��l<)�?�)!6��"�˥��քi��=.���N�V�ۆ_&nxa���v��!���{�iuZ��'x��7=c~c���i� bD��Pá2(ϰ��'���[/������'�4�F��6�NN���`����K��զ\Y�3=�c.kC��p��
tJ�nN����Y�[2�(q4��}��e�\�2��5�r欀�t��������3�B���2r�Ůx-�rJ<�P��넜��@?FA�?���"�+|��~/IiV���@�.�&n�d���v�pN0d�p�;d����D��g�.�e�4rՁ�T�1�k��:|U_�����.�	Em!_��`��W��<қGj�����4qPˊ�Y�N�n(ڪ��O@����Ki���K��Gl�2���"]�vI�rָ�4�ڋ�E�Q�;�=r�j�����
���x꺱���<�Ċ�-\.��Q���~�ۢ[/\[���3؛2��+s�VRs���֑c{��;��+�����X�8��B��ȃq֣��"]�$����%�~��y?3��S�Nb�����T1�0�MV�ݫi�	��n2ݽ�Ȏ�$2���G+.C�_H�}�.������\$�����ӳ���s�4���I�e�6ǆsb�i��	�˝:֡�vv��L	{�<��o�N���l���֝�P�ß�-�biّ�/j�t2BS�zӫ�p�n�0��!H3�YD�u�Y��|���:�½[P��t����#N�������a})�8TT��Sޚ!��@����U�g��W���<&�[��m���5��]^����Q��N�E#����������D���ө�F��(��B������Q�	7�ۘ_# �����r�^B*���~�r/#��Z��۝��F"�B��N���d���bV��5�M��ƀ�ҧ�\��ұ����/�C�7a���?�ذ�u�6��R�N~c64��m6�����$9������.T��u��w�g�U��XݣS��Savvyi�#X�9I���Y]����|�6:����X�yz�M��0��L\�|z��c����?�+-�%���-���5�����o�)e�d�������>�'D ��� p���B��HtO- �b��}����:�����JS�Fdc^)!^L���%#ܧ�������$�f�cr~�4|����?w��DE+�N1���z��z��18���BB>�����٢K\i�T�����
M;�'D�p_M�E��׌;n4>��0SJ��i}�U�P�!�ٽ�����2P������,�0���l�v�>���_�0o�߰��d�XM9�3��C��p���ZL��y���7ͳN�]����mb�z��d�#��6�7���ϥF�?�7鎛�=�<�W%3=`8�C�֟���ؖ��]u���Q-0��_�+-�z��{*e���X1����y�+��0�v��[g���'�Q��]\�.Hlk�ںO��-��B��9�5�E�&N��7��n���E0r�
+��q�pk�f{|-�Fz1� �L&���2wI1�$�C�]�*:S_���1	�cW�
q�ޕ��OG'0�֪���X ҈-����|�<��YI#>��V�rw3Y8��U��Z1�!*���X��ôelD6�*���4ݛ�����j��|�� ذ�H9�B $�a�>d��(��-j�A�E�O(c�K���p�[��\���Pr�f��_u}Ǔ "�xud|-�t�YEe�X!���(�\\D���ӭ���h�2j���Bؒ{ë�ne�_@Fƪ���	���5ҩP�՛�:�eS.Q��<��_��Ȫ'ma
�h� ;6�����%_�{?:���(E?��VX��:j�IV�?a[�|�t$SF�i�9:�t ��+R�p���h��O�N!2E_���B��3�Ԝ���i�a\͙�O���e<�T���a������L��~)u(�I�[+�t؟�7���&����n&F��72�NJ�C���M���&B�����ZZ�76΅�3��m�
�7}3�p�%���8�{c\B�A�
�'��YPAx�K�B�-�X�S����O\�;"FԽ�Ue�h�k9��^@F�Ϩ�ｯ��9߿�G�CL_>��ש�~��[�A��e�z���XL��d1a�,���
8����|�d�֦梑sVl���EK��\��	��ݻ=��T[�u��2��� P�tw���"GQ�1l��],z��Nf:�xqՈi��k����/�ht|W���nVf�~h�]����KJ���ƣ�������
�����-��#B�\z��ӯ���,���9D>
��I5�V���⟬x�]f(T�ۉ�l����vw´XQ�Ȉ�v���<�6���F����Κ�h�0��Ry�y�(ߑ_��凯5�:F�{��/��"gz.��,.�� ��@��!��7>&
�M���*��cA��9�E�U�G����� ~X?%�TZ��e���]�G���[H&'v�m��ț��b>�igB��>(Y�9�Q����U���[>�}y�+g��3�:�e{E(8�3
�$�z'I�6�\��Vl���o �8y��1��{�fu���+���x�D{�����C
�ڽ�#���,�Vُ��5s�Wx�#Z�� �� �\쁋�k���r��?�[�#�%-��6Ms?�?��_�]��6	�����M�9���gcB����0��� �������*g�TSf�Mq��
A}����i���-#��P�-ԅ(���i����+�*'��-W)*�F�����=b�����[��ڐ[�,��N�T*��c�+���s�悎! c&�)i��q�l/:������4հΘ�$�4Sm&���=���YO�������_�68��_#
�q��v����c���6,Gtȥ��W�D���`/�-��ɿ^4����J��M����%����	^�r�KQa��r/�ǒ ����{���7��;����199�E�IЗ'�}�]�	DDw��V�_Aģ( ��2�F�ɔwF�oM>s4mb����}�G˳� ｪ�5C�a�s��u�j�G�c�fL~'1����Lv�հ��·X̜0�
*���_�= ���/�hC�E��F0)D�c�P�eO�U�����eA��;��_����7�r�Yu�����uv�Igv��"{E�l��	��$J�<�Wf�̝�f��{`��n}��}&��i�]�PE�{��hzG>�b��1���MD��7�T���@�e}R�(ˈ�f2�O�����F��]�:P@xR�ON��l7���Եy,�qȖ�	0� �8�����r򭄧:�V�p�|�^��om�Y_1{UX���z�7�>ɷ����D�ƫ��'g���̢����TZ��=���pgD(j��A�Ԡ��\������`컬ݽl���c�:c�|1�V�2�a'l'6Dl4�m����W���P�D��!���[�Q��C�ZɃ�
CJd�l3|R"�L��N9��Y�\;�O�rCH1��i�Wg�	L�Ȍ��R�����"szb�U���%e���%iN)1��' w�,�������Yx���Bjd�7��y
�F�ZS��ÈCbbH,� u4L=K%`�d:_��&Z�{MEd�i��ި��E�3��;O�����y� -��ݛ����̼6%���g`��O��W����p-C�B�r�����b$�(�8S��#<W}�M������@��4�3\�$@:�Td��߹��ۨo�g����]
�'�1:�3R�\�誂6>��B�7�	k�7�#�A��hySV���A��`0���@������T4ށ������Z7k'I��gG���N`Ki�M�D�&)&g�b�R����N?��&V�rx�\1L9=�xyKR������b<[���FTP�P�m�9�l�] `������@k�:�*����zU9e���5њy.�$��w��g��)Q�p;dZ���5ONd�u,+J<��5����� N�4Q��E�T��DNx��k|������]E�/&��kM��"��� #��@2*��	��]�9ut�	Y`�����#���w�a�b�(o�
:D�p
�\H
L6$Ξ��y���:So����ս�ְ��/�ߒ�Z���8��5�!s����o�?m\�]�g��RSj(���ơ_��ol%k��I��~r=90�v�!&����?��i�hOv��]�Z�!/�Q)�k�>d.}�j��B�����?�t��(SoB%;e��/!C>�%a��4�f��q��rBC�llZ"Kk�O�.͋��jG��}G�Z�i�gꅺ�ga�Z5L�,�*�|�}�Z=o��d�?�>w��742�|9pA��K	��S��
`q�8�4E��WQ����/��")�-:*���h>��*�r��#��@*X�+S�9@�����3#&t��Ym��HXlxVHYEB    c397    2030u܂��
p	��_s��`�):,�U� >���~y	��	8�ʔX�R;?���x�����f$u�l���Դ0;ш�nL���> �,u��.�h��(΋�es�b�>C����(l��]��m%/�૵<�s�]��~ô�`� ~}�֪Y"�B~t@#}�1?�X����}}�D�~�ٕ��ͼ�}ˉ;�V*!�Z����;mO�P&�&"^�i0�ǡi�j@V�C���g��ڍ��]�����l��N�t���J�֣�b�BP-5�(m���k�nZʠ�F����ɎO��yj��F\�keOSUCj�B�q��N$�:�a��M�h�W�ohZ��e�	�����$�$�K�r3Z����/��Ʋ)6��;��1{HB��[���H���S��(/&h�����ޜ�}��+{نU�q@��ld�+g��|���j��V�ͯQ?�J!�PGĬ"��g_����t%%�I���G���m[@&�'�����]�(j&/�5��b�����xC�ͭ.203���Vm�@[�>��:�%�l�>.Vm}y��6u��:ks܎��ٻ�drV��n-�KQ��&Qw�\h^��އ> O>R�#�5���{f��5��Mkm3��H�0�/s�*��iY�g��ZȌ2��)��PiM�i瘠���t؄�	�U�r�2~F��� >�˖��GX]<��Ֆ���Fi�����(\ �S��6��$���ɖ��#��Y��E�%d�Z ��d�[oX��{�������L�����O��p:������5�y�ԏ-�Ǭ���
:�@+W�~�8��죤�8oZ�V����yI�*G2����� W����\����OpR7�އ�4���'�ʡ��@�w�䊮��!ľ��%�m6Ջ��#vK�>D$)�+�^ͅ�c���d�< �G_�6��Heb���^��zNvT�8�/G�Q�E�@�������͢��xSbZ�6N��D� Y��"64� �\�mt�-�+��OAF�����6B��祺]���(b���h�8��Y�𘿘+���@|��OYJ�1�D��.���!�5�1y0��X<A3c���e��;�F�ȿ��W"p*I-O���<9ܲ03X����	?�e�')V5rR�n����z��Ƶ}I���ŗt�Ĩ6e&�3�	V�m�7>�M�CzS�@6գͩ�ts�'ב�lE@%�����Z��X�an5�{�[���.Ĳ'�|ɬL�`6�nuo:�E��M����:"4NG׶�5�qKt. �y�řPTxx��q�J�Ӗ6�a� ��v�aL��ƃH�������?"��;"���o���J�RO�A�i��i �P��#�G2�lr.+�U���u�ލqS<�$e�#z�΋��5�r���X'�-d�:��۠���)Xe"��x��9U�X��¸�ȏ�,1�H������E��1��J��}b���e���������cx/��������l��G���X�{��Rd�]+
3�n/|?1ᡨX״S�������&0�>"Aჼd�F�ތ�M46P7\��b��N\�}LsF�ۨ��m5�LE�Jq;�5��o����4����6��� Y���K�'H~�$s���KW[�m�fN n����62��&3d�+�������{�!OQ���㖶2*��.�OG�)�!W���`ŕ���/�J��@�Y�ʡ�J"�Q`���R��8Y�4"Ҟ%�?�21ͪ��f�Z�K�t��uI�T"%���4(�Z@tV�RػB���u���A�E�0颊��Y�#����BKĠz���^`2.#�
���X�.p��	ꆩ*�J�J���@v�s��B��>�_�٢��8����!3�A�S6[�|�!�2��1PS���>=�	=������2����5sO�ѥ܊%\yB�Y�����Lf��+FD�Bg��C���A�<����6�~��V��#��rp�r9��r~f��[�E�@����F��������_f��l䭵B�ŗ�t��vΐ7�3_@�?�T^�_��_�Y���t�U��ân'\��G�&M߷�]�H>��_1����J��tV��ٖ�J��Ρb&Oǀ4��L*Xu�N(0ȫ�Vh�J�F��=;J�i׉��tG�Q����Y��;��9ܠ��G�r�T|V{��C�S޾��y
u��ٯvAG��ݛ�ҌYl�B<��_�[�FB�Uq �+)�|�.�U��p�Ԯ\"�n$u�X���H�'�W�`(E���(���Dݏe�@��n��q4��X\lvo�NʑXc��i�o>6��d:�����3gD!'A9�ccv��NbS�=�J�<��̋g� ����k��Q�EOL� �O�6�S�-� �y��L�
kc��rG��){Mx��Tܽ��M=�r�P�����������j*�V\��U�/��ٰ5@U����H	G���plL�I�^3�M�d�tϞ��"7�T��K�����G0���� �{���Z\��^�[�����x[�)���@n��΢8xн�\��/(Z)��Mn.t����G�9C0���O�=�]����|�BQtL�i��]2�H�P�Iw�*p������nV"��i�W��q |�?1^|�y�ڞ����*�gg��gg�Lwt{�,�䊬������7�Ǜd�ekSwo�>ėb\������0���LX�Z�A�^n�,�r�2��Ww L��m�f�2�ı� E�羵a�@� ���0�Cu(�46钖��β��E1t�F1��`��V�V%�A�p UDp�d��^�X<�X�袁g��;l<mq� Z
��D�Dsֶ���[���ykk��dO�)J��-gSDE�����, ���`ϖ�����e^�&��� ��,��v�]�����w���D�-�6�ݎs���k)�`�����a�k�P�EA>�I)O$�{����TzY����_�}2�r�;v�� 7w�P�Ǵ�귆�R��vk���q$���9�T��|�0id D�E�E7@w����k.���4XV� }��>X�~khyL��m�}�z�>����ʒx�"��v�\X��a����و3�S�{:��~(��z��f���gq�2st�y��4p���O|J��� |�N}���
L��A.d�")���Ha�o=Pg|t���$������?��PIS��;�?^�hDn|e0�N�� &�\#��I�d��� �E�/?�5	�O-�T?vb�.f�)A6���0�C� 1��`��U<��i��t	�Ӗ[f^��(�n=���[�N�x��a�����$�"�C�,���\γYFG;���8��dB� �>k�}b�}�H�1�ඎ6��:`MB6;�W�̛��_���_ �5��tAj�����jsCz��(*��S�8���Bh�ݪ���ö�	�$q�#�D���$ +P\�(�7Fc� �"�Ht�ݐ�{��z���w�o:�u3y��еe��v�F���򶺆>�U�J�\Ou�1��I�����u�
�r�G��%�0����q�u�7�@���ن��cB��f ��ۍĹ*K>D��j �ןSP�-Cݴ��Bb�<����	0�Ϸ�j���������{&<��4�l���I�i�X�A$�C�e�bh�W� �%G0塪$��F��<8��҄�bf��e������k,��q�2�%&o)���$�li���9�PT�$e퍥W�:��"�?�/1����Mc�Kx�G_�>6�1��"p^�M:1�,8��z�z8,��	�������̳����B
��X%b�ƫ�e���p5M����	묛����hE��x���*��y\��^z�0Ů���|qV�o.���:¤�alXtL*#�����f7��/�&��^��]����Jn��E(���_P���=Uo������
Kl���� m�p�mE�8�Z
��#��
�B��h��I';
"�'�H��CN:2y�c�7?����Ic~'�GA�J���35�	����b~M�r�f��]�I�	J�`L5�ZyN�M��GF���f�ZcT��`��x�u�/Bu���&����C>�utH�\"�p����ڵ��[�%��!k�Lm<365�x�%�\�m���G��QC0�u?���p˷s�.G��Po蔢��Cw�U�E!}�X��c��γs+6|� //g���\eX��.d&���^D�YҥB�kÕ����?�N�`9v�$Oph����0g��} "V���j�)�t0&TA&'�cs���I�^��j.Ӻ��\�S$�,����fr��&�B>'���$]�CĈ�ϼ�F��X=Q�FG^c�9qN�g��$�h���h37f7�4��V��l�P�fJ���j3?wG�q��F�_\�KL w,�����BhN$�UMA�-�Ңuf�Z�K�������l�๡��oDlO�_X�?�ڎ;NΞ¶����y_����5ď��X���|�ΆxO�e&��,e�	d�]�]0q�+��}|V�^#�2@�a��#������M�NQ�t���'Nd���|���m�O=T��[}ϳJ�f8ræ��j�3[���{
,r��kRC���/�u��n��m!.��"L��=��
~b*,��1�� �o�E|�a)���˻���Xh�����oO&ğ��c��!"��~n�B}�	��A�Me��Fr���mR<�j�+%Nz<�>q�\@l�ۛ9��N�3l+ay��8�h� ��dK�@T�}��=�	M���,���q��f�+ ��6J��/f5�>p�X�.Ok�LV;��ǽ���=�� L@��tw������ԇ�_�|`�[���RW�ѹ���H]����{�<fa���%�j;��f�b������Ef�R���c��˸Ѓ»/32��tE�tP�W�u%&B����_NL���^�������$���u�,#�M�V.]6����x��*M:�Zfx	l3�B8�|�b�Ǖ�|0 ���Ð�����%�g��y-�~�-���s?Ρ�c��˄���`[£f͗�dx2����n�Q	Q{W�/�x��4����TEW�K>��N=oz�Ry0ЭU
W+H膠.*����䯾�M��ǭ���6o~g�Z@Ԏ��x@�w�B4���.�򠼻��7������{"�72�ĄS׉��8���њ��O�����3�x13�n׿�^};��W�^�\�Mx���Yw� &��h��|��	RE7A�@}�B5��bk �z�;S��.Q��R���8`u����TA�^U�/����&����5����6�~�5z�T9%��l���X�P�6�GzM]t�-��X���J%�v����ʰ &E叽]�׼���˔EO��6��?@4��U�s�/�` ���J ���7#Yh��\uav*l�+y���|n��]/@�K�����MAH�R%�Q�ӏu�,����Q�M��x���5�_=E��S��Mb�x�\G�+%*"��^n���"�qy��~t�$��\Ü�b�K�s�b�o&-����5>�][��gB�@㉟c��\I�kY�H�`1f'�-��꿻��nq�3���60f�S/�t�]�|HD���\�c괶��FE��������h�*�H8]M4m8
���aպl������f��C �h|O� �D�N�{Of���4@t�b>3�N�J��I�+����:���\d�!v�����,-X 6y����dF���?����Ȼ�������3��+�͆,�M�{I�=Q�|�?�%?�X�1�m�1:��l��:�2��kԠ���l�¸E�V��H�tbo�v�Q�ק�f�{��:�1�<���m%)��h�u�~ݕ��hZz���v�'�fQ�t �Xwp�4��LU��"l���nV�~�7�0X�I|U��_%��q��/�D<�w�Tw�,�J&,p|�E�g��z�3�����C~��n������t�S�{
ϭ�D�e�e�f�?$��&:�$/-9%�/�>�r:J��wO�����!�I���5�66k���G�@{���ּ��]G�IS�Ca�����xZ-O5�p��D)���L>��/�㼫�V-��Т�M�@D�b�=���懵8��s����K��:�|�v�{A��Y�93���=r������Cze�YkͶΆ0���taO�ihƠ����D`߯�E�[>��H���(�Uf�Pj�N��_��}�Tүik��&�NwҶ�x��A�㇁?h�B���T��e����N�,R�����f����9���,��p@��*�S��'�{x+��<����G�>F�'n}��K��݋w��"h'r�ǎ	m�؇��TғOgUO�x��j��)j��B���!'�)�@��rtκ~ ��Cp[�e�A��RA�7�7�m��˞��u/B�¾�e���$Z��ܥîk��{�w<q�3��D>�����t��1_���rѱ/6�����Fb�wN�CŤ�	6�x��9R�T��˨�O齈�X�[\u��Gj1��X�gX�4>1�<4�Np���9W�����I�x��D��6�p0�:x�2!����l�r�� b^�E8P*T-��[%����^}����9�N�0��-'}!��@���rJ��ˈ�	ś�h�%�l�;�cT�$�Y��qŵ��y�tʺ�C/v��z�t����{{��i~��{�ifR9-����e{s����Qq��m��9X��p��	��=��bF-�tp���jJ&y�>s��	W���Ԗ�YJ��O"���Z�X4v�d�r�-T��&e����Ƥ� �""�2e�l!"��ðjі�l�{��f����Qϙ8��Zu&x,@\�"N�|f�	�����#�&Q�b8K�h'�&2�m�<��&��VYi�I��6��	�Z�{�|&�=5���	$�{�}9���[�
������gXZ���{Ci�bCۉX#d|>n�uWj���X��"i�9���sei��~����6�����ň�����U�ȣ�zt���f.%(��b��#g�jI���+��:��)�if�X�g��_��5{;�FA�Z���p���)c�Ff	�#�Pn�f��'��[��TxMJ���;`���)��3Uh
!�E������S�ru����c�,zHL���tN-^D�l�
˰J��K��u�A���
������B$��,�d��A��2�����;�sL����Q;�@��ħC����λ!����.�r��t��)o�Kü*V����j�!��fz�d@���NlEɾGvF��Q���|�mO�yYq��B�u�u�o�����E��K��}*$W��B���w,�Jg�kr�fj�������G��<'����Y�%#I�<�ϼ��L��b�B�?�ò�/fĿ%#�-ذ"X�B��	}{�rX�.OO�#��T� �O�OA��	�v��z�Ê�sg�c��L�($��.8�B�C�+�V�^XqC�ȝo���V'�w4�(�^ܥraID����� �~�t��!�␴B�7@����[#0$.�C�a!�P@Ē�LzJ���O���'QI��bh��e(��}Yx� ���BJ�$���.Dc����Ai��+�L���(�Gxc�)�4U򑴂���㼭�ZE�V~��cq���g;�W&�|]�-N�-��Y�m��gد<��ٷE}ka��e���hI$Wo��,���R���$�7G|+	*"�����lZ�ʈ���R6�dӭmN+c����I�z���q����Gk!�fH�R�S�Ѻ��P��8�X}o�<�Tj�WI��8�-z/V3U�hcz*��7h�_p&�F>��9�X��12?�As|��'L�v3F4�7��|�#t�R��� #�R�-�H�'T$������D�m��{ra�0���_ �dy#�`��}w�\~E��n)�s0���:�[�!��W����T)BU#����8��
����!8��x��RK�������oIT~�����?_B�2��yV{��\nZ,�p�#ŨǴP
�?`&X��#�k�)�fG  �|�"�{Q�<lޱ�c���(��J���5��ye��Ի�u�