XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ü�r������YM��l�RV�Q�2K��N�OZ
��V^k��e��+�:�����B�gp�LK�L&�-�ٛPoG�d�=E��@�qJ��+��3�f.ـhs��sxiU�?@�ܬ|!�8��wJ���3��0�����nD���L�2��&� ����_��{�Hk����\�ԙi��� �V����m�l{o���GA%z���Y�݌©�)�t�K�0�Q����n���MU��vA�J-�ʡ��m�{�����$"z��Q�O}�t�g�t4���2�Sl�#f�[������X��ʮ6�UGv_,��b����j���ؽ�(c����1t�<S�(͙���K��hơ��0�,�#^<�aI4Ǘ�yg�?��1��?qgs׀Q煩�.+�,��8L`j�Y����^�	I2E����M�œT9�Ec�O�hE�'$`C]u� �fM>�ƅ���.Nq��.��d%KE/L1�%�@�?eɴ��!�"X"(		q�����M�;$����9���w$�.ܭF�;c'���fsc�ZŤ{�6 �S�#�%��T?�0D�c]�f=4�Q�l�Zk��M��V+2z@��ɇ��M{�@�@l�.F
�7�.cd�d��-⚼3�XX��P�|�� "�Vv��� �mf�}�;p��*����󞁡�i[�([����=��W��)pn�Ojۢ�-��r�����g(�#D[²M�1��Ha/d&�'�����ʀ��tA�>"���f�L�=�&��؏�=�s����Du�XlxVHYEB    7a7e    1af0m8�wVR�^�}K��/kc���I�ɿ(��%?G���i�+'K�ܕ��TTr���v�)��>�� �G��< ����/�K��}(p~/��T\�Ii�/4h{����gj��<=��(��ir  ?lQgv9V�?�L>q3���Y��0EP�:�!Ju2Uc��{ʕ�jC���jDQ���y�H�D�Nv�p,�Y֠��̖ >SR�KPh]2�������H�1=p��s4�Wғ�³.�E�-+��T_�˨��'J�Ѯ
���/�5�� �k��J��)�J�0� ȫA�HM��Y� ��?X��hC�V�N���K������k����M� ��̄)e��Ll�>�uk�6f�%+A2"ˏ��ę!�|�������U��1���Nn����������$O��WDԥ#����s�	�g�~�w��V�~�IF����{���Vݔ/.A�56��_�bxG�n����U-����>؊��Q?� ��Y7C�ͷ�%m��K�n1��y���exZps�!Bc�L��T\S�ʋ|,���<�G�V�ў�I��Kb�M���X�Ӈw���7�ҵ@@Q��[�rѢݧH<|I{2U<�uD
&<.�3�?����o�*���2��qw���V�~���hk�.��j���M�n?,��c]�e͋O���K-��eZ�gO�*[iך�����md��}�eK���.�ZG��ǧ��k�bQ _�����q�y����_e�n��.{�Ka�s>^a��Kfx�ݬ��7.(�Ng�M_v8�b0�Ve������@�3l�f�[��1���qP���j�7���t#ܓѬ���_\˻�aE�t���%�-P���:�e��ںɐ�L��wp����G���cdcwĬ;DYA6�ɤ�1�D?�h��Az�c�H�����T�-�̠���`(�Z�L#��{�3Q��VR}��/���x����w�/�P@j�F��I?ӓ���E��{�?�7�*�*?�4x�es�Nn<�*uc�do�#��Nt��w��۪]2�L��h���G�!������)�H+I����o��T�L����(��e�E���?��ƎQ`j���?y`��d[��O�3�� �-5znc�K\zV{�b��VS�������m|b��'"L5+�L ��xqu��p�8�u��m��ej�z%��E�ݡ���E���;}z�K� (�����X:�Wj퓝�Z�ٞ��߁{.��)d��;:��(fفv��}=]{P�1ӑ�a?�Xh�u�@ֳ:���j$d��"�G���a`]���[?���@�C|��8�L�y��ձ��R��M�$#y��n��&�%��u�9��EHvX��:7x�đ�L�/�'S�SxԵIn�ڕcQK����{�Vc$�>��7lr���＃=(�=5�T�]-^�<�x����o�s��O��U�-��ܑ�L����k��bf:Cj�%+�)rih���D{L�t�X,Z�8�u�^TDm��0�{a&����w��)ڮ>��K��=.�f��Ծ�C:s�^E�f��7�x;=������	�K���l۾�>}�J���	�}ޓ��}ʅ����qS����;|��,<6�����:����d �y�������z����L��W楘@No3��Σ�U���c	t>��� ^�݀��/�Ьi=�AobԜ���XiY,칣X�X�~��!��Z}��i��D��t����K�>�&�Q�9�h�-A� �άs��I�$	t!�`�F�Q����� Q�m~Ҏ���ܠ3�X-��F��%�;�3:���حniP�AV���ACv�^�T�K����~����1a5!f��t����r��퓅�q\#�����7�nO&{������y��P*`9���q��)@@B`��c�R*� 9�N�tT�#5��n�=)��o��9�ڪ;����v�մp��>��ٗz��t������[����b��0�U.���іo���s�:��Ժ�c�L}כ7�P�|�Y��� ��%H��J����?����ͥUN�����|V\�X�6�$�[$��Ì*t���յ��Z���(WT�5��ߨ3U�L�Ú�7��M3J��/t°B��'O�*M�v�{뮚Ct�۹�K���>�A����(��2�nҨ�c���Z��K��E��"�E%]���e� �6�m#���m���G`�;�A�<L���8���U-�?�ob�`����үw/*�HX�&4s̿��Ƅ+��m�ς����czTzð�J �wR�i� ��O�{�l��υ�������Tu�h��K>_���8�t-S
ޖ��5����*��;��=���s{qHY'�_�JKsn<fN�T4�$ʴBr8V�A27�a��tk:8ds�c@�z�!]�����.��=[�h��ojM*Q?�=O�[��(A�m��2ďfS����$��@H#�	�{�VLv��T����x���@ȓѷfg$��O�E4:�H[&��z|~]��kXLs~I\I�>#���R�}r~�4�EEG"R��zĳHX1@`��)���B�Ub���	��V���+>�6�cEbE��}�]�3��ق?&�W�1.w�&�I�^B-)R]�oL*L��
T�(�]��*�Cj�-�ͅ6��=�.?�Q�ElE����xf�@�J�8�G=��J'���.��� �_�|P��_K�������
?(��>�v�*w�|�F��}�����ƃ�kiS�LDϘtyrXKVþCh[�2
���+:GC���_��x�޳_.r�T�Ϯ���d�,k�&H�(3BF�.C.�မ,�^+f{;H�����G�Sp��>���|�8��Y�-����ܺ�F�PS�C�����5���Ι{��hծ�}k���@�g?h�&����Q1�"�iT�6���c�$=h��(�O���m�p���W%sD7M2$�rT �l��V�I�@���2�5��Ρ!�"J�%_�C�1Ǟ10#59ߚv�
b��s`���	�P���V�*�6in�h#-mg�IN��D��?�2�l� �M@A�`b!q��hd�K�'����9)���~���:�o��eR�E�2�C,HpW����~va�G�7�r��� _���'�(,uֽ���� ��9ڦݜ{ �Y�m}�uM:���q�z��Ѕ�9�\�2g��$0�������8����ժ�����"Q�/8�����\ ����Yd�7췁����c��60�PNw����y͡K������^L~J�v^bV�MF����pU����V��߿���0�TWT*�*cK��%�=1�m���98f��2����PK�h��AP�u7���z*�:>!u_�7�c��#}��V�Rfk��f��G?��r���Q�r�v�+���3�}P��ܶI��`M�]j�3����Z�ˢ`h?�����liR"�w���Zx����;���&���y��� J�0���)3���3�,tJ�'j]���-"�7K���"��$�f��q�\�Ts��M@�ⴭ�d�����
{y�XĔ�F�-r���u�(�,�1���0z>R�L1O�{\�"��#Z0֪JUW"�p+I���~Qq�#����oq�)0�����Ύh!J&��'^|Ҝ@��!#]�,�f��g[4� oƯ�'��(�>f��=�[ M�,y���(it�4ڲ����%WuR��7�n�uH�7,�t�6��,���8%+з0��9VØ�q�lܶ��.�k坚%���BD7��!.�E#'z�^�Z�ݽ
)�e 0t@�n_��[�9AhkZЙ��yf�9���E-چ�6�O2D:��s�yz��+'p���%v��G;b��w�I(���?ׁ�,���f�X�$Z�	<��M�2ֲ`�WOF�[��B�z�l'�����Q��j8n\ގ��A hd�B��P�*��Q��?�i!�Sj�
2w��A����-'o��� I��ZW"n=�z�}�ww���&�3���اG�q[,B���q�����-�C���3�J�X�6##�Ei�Dt3��{�@���EX�"�'�@;�Po<����cF=~�����7��q^0�6-R��e,��İ�5~Z�V�K���_�+���,D�h�{~V: �_�M�Ĕ&g�ˬĆe7QUvda!�c��b��Ҙ:?�	�a5�]@�B�pP�#g.u1�Y(|��+B��0 W:��@8#��EX���nS��!�R)~O�q�p��Y�H��Zo)m�_[^p��N�0��z�Y�h���ƒm�Qo��yD�-�վ��Y���nl��W����X���!Z4��@?�N9����6�0gf��Y�e,���^���d�@s�6�0�z�n_�S���0B',ܛ���sQ�:-�ǳ�795m�$�%�4�Sfh��_�=D�i>����4ݕw&	�Tus����EO���=�+�q��U��> ģ�O�FG�����+���GY��Gb���ފ�j���˥.����C�-~e�8���k�H��SɃۀ��ջ��9!���>��2x������8:Gqo��ݩ��7'[:,�ͨ��Y���)�cQĜ.}��+��e��U��7�X��X���60��&��u�,�� ���07�h�'c���R�!OW5@��'�v�@:�W
J�~����ꀊ�^ �=n0;��(�ZV��}�`��o����*�#�I�G��#�p�ؕc����X�[_�2�=v\\P5yJ�y�q�g�Ȍ��
V��kv��c�ק��4G�i��	���b��D�[EQ��X���m���������_�_�X�94-ޞ[M�L���k7�f�~s�9�*]�X�EF����#ӛVR��x�C�Ɠcƹ��;��!��A�0�}���V�q�>����R��cF�p�\S.���z݈����~�x8�I!�D���pB0�xЙ����W��L�R>�A���{�u3��W1Бgr���b���5����
ι����9��m�Ѐ�`X!r��v�p7soCMZ=��0���;�dY\b�=ͬ��u�X4Ut)��K3:S]���\
 ѐ�[���L�
��.�J��Y"#��˒��qt*���q����߳���vފ.Ţ�4�V�''�a�A?�!�t�k�����2�/��|�n�gC�ׯ�T�ܘ�� �K߄F5ɥ�JY{�u�w��9pYb�Z0��[�ޙWP�� �9�
Z X(T�K������;o�s�T��3lNG#\���6hkr/�w5y���+Ba�1җ�t7)_��x�6��EXNP��6��?����~�����g�j�R�"Khjé�����@K�%ڞ�|�����5���*�0?��h��M�)`zh�eɢ1\3c�.+��/b]�\���o�r�"=Qr9�V,j8���K�_��+��T�V!��uM�%7�?��&����x�qU~������a�N�н-�_E�o{��xwR�2���7���?�Z�C�{�z����O ��������(?DZ; ��zВ^��4\����'뤅O{0�7���i⪛yJϕ�x��t�E�l�����U-5V��Qv.=����iD���&���9�Ո�z`a��"ݔ<ez�>�Ʈ�1ʚ�φ �w~�6�,���xZP���kh��H{�p�ן�/����K����_�X��g��Z
��(��XtW
_��P�:��։I��c�R� th�r�f�ؗ]�z���Ӡ��&�/�w�O�w2�Y�
q+�&��,t��&^�	�'���Z�h��q�©�I�%�3��w�)jI�R7��<��gKFk��*ٚ(���9���|T���a��!ɳ�����Ui�}Na{ݷV�.\	�!�EM	�'���`�S#��|�Ȥ�"�����U��u~=�5C��^D��y����@p�e~ٿO(z��'Čۡr3��U��;���8B���_,� A�XSY�d�;�~���HD�𪴄3E]���XÛ�
 潾$`�^��UU�dk����A�]��UvՀ)^�P��Щ��}�p�;�/���]�Lg8��z��`����0,�1�!�y��M���/6��Lc�UҌCWX�r�a�j=�_�Ӛ`	�1y�'$��OH�3�� �.EnaQM��Q��IpH3�J���dM7��0�_s�~�����d*��D�[)�B�s#�EL�[t(��{!�������#C�͸�MP0Q���M�8"��n��@K���r�˛���Y�+MV�Q����(!	�n���2ls�0����F�:�I\�B=��5o �-��䙝��z(�4�G}�Tv3������i�M��xEjY�Ҕ����%�䰭t�Eʰ��E�BA�kԱ�(&�J�ş7�F$j��']��^{��Sޑ�_���#��������|�͓���h�!)|M��K����0F�ãu�N�&�/��HF��d�q�/|Q	}�=?�d�� �I�=ԫK��f�G=1j�:��}��4S�~�w��Z����Cz���
�$��F��K5�ǿ����"^K����d�"y��{�3L^,�)�2m!0�ȍ�Moc�ФAS���xx44�`�)�4������?��B��m��J6�W�Լ�,}8�A�h�m�o����_�8�~4U_Ch���L�,X�	��^���?���Ҕ��d�s��~-��h�r2��1h�d>�r�t_1��.>�}��d1"��x�V��زth_Yd��<ju���XM����C-��+�� '��M�&�(L6@����وC��lm��Z�Ap�M8�K�dp5�����o���iFO