XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����_�Kq����F����I����X���Y���OYS�o�F>gE�s�^S�л({_���:��O��p��f!Z��߶�6�����{?�=0�G�XW�p#Gc�����9�Ԋq �/q�,�*���= '��͗�{x\1l;��>Bi#���������z���h*S;��f�Q��C��<99_�}ՃɼK�����H�gH#l��M�_����٘��N�OŜsi���9�nf�����-��yw�����꧀lf�m�!. C[���s;�7U�vC\�&�vV@ �#*�u	���}d2y�l+_炎��YW�p��4�ט�sk������f�ٍ����en"�w).��t��wY�A�L�+R�����.V}U�À�6�W���v�ɓ?nu�B@�j�Z���*�'"V�ݍY43_�S�=(�Uͩ�S��=���zB�pv62�s7�B%w[=�˴(]�b�1�Wx��,�W�*_4����B��q��9����IA�z�ر�ҵ��93�C(��7�����Vq8F{�+�w�iub~����ц��L���+fV1[�<�o-�4�7���[Ѝ����0� ~�������3�T�!�]Z��6�f4��/\/�깍Г^��F�L��k�㗢����f����U��e/)zmHs7Y���ߤ���
b���И�y�����m[]=��� ��A�����%0�n9�,n/����!��c�<���*l/�4u �4k��՚�U=�XlxVHYEB    6ff5    1760$��u/@j�F5}v;] �wY�멭�p�(�r�(!h��K�`E��ez�V���FaF��q�|Q�2�ʶ�NL*�q���ȣ�s�E�J�g�ԑ!R�����l=v��H�]냝���e������֫&x3�����F�G���9Ӭ\���,�2�J��L�/,=�O=��$�?�s��K�a�}�g�#��Tr\Y]"�q<+�s,�zܰIv{'���V���:ԚF�3�vu����#)��N�2~ͱiR��vK�ŭzD�ʐ���R�#+��
������A��,�Ѐ�\��Q�U��g����B�E������]��E�o^���!�@�ڙ���1l2�)g��[D
��1���u�� ���*�O�s#�6-@�d���n��*�,�v'�ZQ��:�q�����m��2C��M�H�D�4��Si��wlɘO���$��V�k4�1�S?��N�i�:��G+2��ٸ��H8�
�!F�)B*��Pvbg'�$��'�'�;m�z��F��U�;����.Y�Wi�;�)xXބ�A���m���߽��Ԫ�.�,Ԃ���$�luqO�=��pL@��!|���&� IS)��Х�퀑�8&8�>h+���ps(��Rf�<{��/�4���yʶddh�Qf{��ߠ>Z�����Td�\#�E.'xq��R�DlO���m�hw���! �Ǟm�Իץ���R��ps��gcn#l\u���k/4��9i�:��-'D���(y�
�#$�����9Ͱ���tK���12���<�柄]:u�����H��3f����ͫL���5��vI.���Z��Ѧ~�ã�U{�YL^�_-�:`�T���$������~�`��*4�d����􉗶�h'��i��3Al��{CE���y"�a�|Lr[S��q���h�Aଫu��YW��{��3G��3m^���_A�6UٞS/4.7g�`�<T��}T?��ps�dh��ۈ������wq�Fp�������M����d�c�]l�2��Z��I���箞�
8����cA�%19j�Ա���Lc���Q�l� �������O^�BH�Y/a��%��2��Z�%��?c��^��'4g;�z�&Bԩ��~�=�����~�����o��z�{ϣ��%* ����U��
�A�xUݥH�H\����$��xiR�)�!�.
�TG0��(o_D�y�+�f.�؍�2院���z���$wl �qJ�H�X#�6�T}{RiN��5(�jO=�L�hò�W_��0�����s=��s�z�F��{��V�(�1:"�L�q���ɮ�*�_Qƞ�����Zd�������q̐1�}.h$��]��3W�=u����;'�B�����S ��c�*1�Yo:��g���<_��S�F;E�
�=l$WX��N|��?2����b?��H��q�(`��X�e	�$�A��]c��1�n�}	�~Bb���4���]�X�'xq�W{��6��
����6iL���A��x�$(wf�|�U{鱲F����p����- {����+�P,�Ҹ��N�$wA�F
�����|�a�ʷ���V4�,vZ�:����t&H-��l93c6/6!t��a,�_9��m		Q�\q�Ԗ�����:�P���P�4-r� F���Q2bC&�wY����9��E󛙇�]S�Ӭn��N��E�BV7e?zs��(�Ϸ�>��;��t/�L�)N�?��i�a���g���[���!?8�<sJs+� 9���������	1;����m]:,^�JTB��u����$e�7�Q뱒��*�D��SA��>�-�Ϯ��4�m#ϑ�Fv�S��cWc�sUT���!IJތ�
�H_�d���r���o瘍�^�#��u��5�e��^�-��h��#�w�kʣ�M�S��p�l �Z�{}�Zx��v0yM���a9�3��f�hj��� ��x���%��/���4�M��3�m�,��S{�il�fP�Z1	�L��++�@��K�������	h��Vy0m��`m�,����w�c/�Ź��_~��Tnn����_�'w'J��a����,�Z���a˼r9cI_P�q�Xg�[�ƈb@�m�a&�{/Ѵ�I�61�jh�V�Ӫwǖ��aJ�ʍ���[="]�"�2G}Ѹ]0�G��#�,W�)AJ�~�;/�*��$�fs����y�xzO��{(������W���X,g4�@ܬ��J��V�?��PcJ��f�u��!\��~d��oތ\��<.�c�Wq�t:�4�䗟�g'u�;�s��4��%��Ƿ��v?AXo�3Ȏ��1��:�,d�SM�Ȥ�5�j���^V�Z�)�{��)���I�?m����{t��g���-�)m���A{���!��aQ�Q��AM��-1�H<�D�H@�NM���d�'0v?Og�!��+�¥��b�����:d@./5�ęP��]a�5�tR��N�1�`#����D�1�jS��R���{mdG}&q�{֥_�1��|3�↬���y��e������{`���}�*������!��G����ȷV/I��{9͑�s!��h�7��L�����/��ڧ��"���cvH|��$(�̴,�믯���hM��,$�YE��#� ���X��ѧSr��'A�zl�׶�Z��x8r7/)��,<����lc��f�5as@�GCi� ��&#����p��I�ro0�@�B`O".�)��聆��K�ChΘ���م�	&2�t���é�dD2M���5/y��R�NOg�yl��^�kXl�\;�{�%/1�BG�b&T�.�K�f��y��H;1��>���H]��3��3��s#j�j��$���j�T/f)�g�?���h���3��Doу�z�U�<I1+�H��M�W2Ag��XJ�E�� ����g�ݦdҜ�ο�u��	�B��
�Ś�4�3�������2
� \\�.X[��^��-ҏ�A�h�#��2�����2��͎^V�m��NW���1`�Nu�{W�ΪՌD/cK��AoOSMqu����$^2�C5�"�(3��k��1K��½֬�y���%���3���5=zľ�F7�h��둰����M�)�G��T��>��%>�^��#>.JX�nbԲUsS�P,�F�~Q�,��M.�(.��Uo�Cm=*�K�<�_¼�\v��?�_������Y(��_T5̼����B�6�ݿ6��� t���:���J�fA��}��~K$QԶ��"��^��B`_�Ats�F����.s��IS��kE�T2�f_Ȧ�L��p9b*}�Q7`��4J4^��z�6i�\2��A��9x��p���'�2PA�,��#꫶��_�:����$W�ΉYCQ �yO7�v�U�R��
w�
ս���aN�HLh��g?L�J�K{E�g;�l���	b�
0��~Q�JX.4��q�e�/��!�5ܘ�J�_5>̭�͢�Y���Z��4���~Y��ૻ�N�t�FF��YS�
�3�
!:��P��|� ����N ��bV�IvF�pY���g��r�b֧���_�W�C�E�JK� �_:E����1!�V��?�pH%�������*�%R�zyV��O��)C�1ծZ�bKu}���S�/A����x��<�)N#�o�ԋa`�5	Ɇ5���J6�0d����nh9����VXY͂����i2����剥��|=�$���i��.��<C|)�#��Q_Zz����8��Ӳ6נ
JoV�׀�7�"c��|+��9�������'G�%���$�!�K�v��(Ә]���Db��9����&ulp��� ������&	>ۭ�:��2D����7�Kϸ����K�hR�L2�W�jַYM6���Z���%"&�ڴW�i����?t?��.[9
���TT��`D��J��)��
�	�oh�TDV�^���i�n�ä�a���p� E�,]j13�-��י�@w��hQ���JQ�m�Lf344"amq�
ۗ�i��_;x�^��}�#A�`�e�~�v�X��=���\y�yy&��Y�_I�հm��O�+[&���2l�Pn;�G9#���RD�8�����y�n��Gy-�OK��[�@�~��vȾ�y]4�����!|���̶�,	��7I�}�ŀ�碨ß���>ڮ�Io@rX2J�4؀�wޜm˞�	b���1Z�w�/P1�T7c!e��AG?�y �`��+M	t�&ףza��N��a�(�jxIxҾ��%fø��bw:̌��Cȧ@�x񅁞b�岷C�o�<������J�.�q�p�:!E�����;4����c��+!օ��wH��٨���D�
,�dh1�:I󙖡��5#v�9�v�	K#�ܥ� *>�h��A����︟�IB4�� a�,��x��ϴVwc*��T�ي�!F�Z����?^sҨ�7!%�6�h����*�}�$[�,S$R�}SϿ�C5��b:x��J� b�;�97y�yP0W�_�?��J4j[m��'��Ly����)�/��L��@�2A�"מ܅tޢ�"�S��#������B1�n��gk��P��7OX<���Օ��w��WDɤ�3����u��fq�L֠i݀����M�&��stbK[�"0�p,�)X�q`�88m��)��!L-����	1w�����V	Gx���&���r�*ܭ�#O{��Jp�};��}�顪��o"��C&3*��w��x�>r�MP���O�%;J8��ǧo�3_�sL`I̚�̆�:Ӕ>	�?d��r���n����I�TWJ�nֵ�x�ԩ��,���,˱t�i
�Mf�_�m�$�qW���jR��D��C�8�����#� �uD�)�El���i~xg�!Kh=#Ҁ"�^��3� %Ӷvl�?=Z�<`�j��EE*��X�y�>vw�I�����2)'OLt��	�r|�z�j�Cw;��x��uuj,gQd�GͮǵF$��[I���ND��F(Ǔ��	}��^����y-=�Y��է)����}+@�� �+z%���y�酥tG\1��y���ô�r�6#��NFܴ&|(I���G���g���_-HX�c	�VNK��/Sj�'����#�֨��J��2�(RZn�p�Ic���/a L���=��L��-̢�kKD��e�?h!�Mvy��6��_x?��8O��QC&#�'�!W���G<>i6�Od��Ϥ��~���ݛ��!�����T��-�Hb�pJ&2FE>���\?�A�^��xt���L��CX@�a���-�e	ӊ��o�d��`�)��~�+�i2c��l� �"��f�D$�#_��v�ߦ嘿U�!��u���QR�{�t-j3�{��rQ�*i �Ir�
�p	��I��������.?#>��Ϝ�dI�L~"��������i2:�2�j��Ģ�A$X�it��ɕ�K���.H��F��$��X������MQ�������H���Sl5X��&y(��N�箏�7w|	,��cA7M��n�=�Sn(� 2�����5A?��$5�YZ��6m��V�\zA4D��]�/:�2��tf9�]�У�.K��,G.q��*κ�Ebj�3�-r4��S�4
��6�!JF�ܴ5���t�N�4��xEF���?ťrv�7s���*I�-�����H>�e��+T�����6���5��s����>R�5n�a+1����)2��g����W ə0\�1z7��fw&W���"d�r$�'&���(PE��sK��e�Ջ�����$:�J@P�U�f-�j�%W�'_��x���1�H����U������%(qL'�����