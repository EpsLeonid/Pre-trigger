XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:\:��}]����u��g_:(Ҕ�8�4{�������xn��q��`[rn�b/#�F*鞫�Q'���@��@��/#�X+�"V����x�˸B,�0#����^��[�]mt��Qf������f=P)gzBQ�m^���t�=�q�K^�-K�E�Ts�W��e�'��+���[�Y�;�kG=���"-4Ӓ��u�e��K�$��A�1��f��i̹B�׬W��r�����:͖�Oj�L����s��4��>�8�o���\ ���$9�v���ﰨ�]�v�9]~6���5�\���S9��2|�O�Y���)y����$֕(S�S�v��Ir��z���{��-��.����f7L��5�fۮ<  2wH>����Q���<�����J�qC^��>�����ڲ���~y���#c*nT
ܺ�L�����Ch�������̕�2���?ꁌ�qe�NK��!�XI���/����a���� ?"�7��K�V Y��^�R��/a���hRQ�S����4A��/�_K�;de�j$9!�4�&��9kF=��Rϔ�%jI�o����ʣ�R9zf�+9|�	����)"�X�R�k%�nJC����7^�物�ޮ�� u_��!���n��Uw<�%@�,��$�-�����6v��P��.���G�l�����#��<�aA� �|V5�o,��p��Q>��K+��\��"�XE{�5��CR���l�H�k��0r%�ƴ�}GXo���z�nӂ�LXlxVHYEB    18fe     880��٢��?�S��uS�i^��$�^؇� 3�c"9�j�\��>|�d�"�5��)����� �|$�s�=-��9�\oR�_��H����F��Ms��Ir�����k��1b�J�X�`�r��N���u�M�Z��5�4���<�i][�-�%��rUS�=�\,��9��F�����5���=���2o� �
���,Dq�Ee���q=`du�x��_�2�����q6Ovs|���.<���3��NS�{}t(��Q;��`���������?�V}z�gQ��=uBPDl�Y�69U���N�g����';�('�{�v+.��֙����W�=ᾸG��ɪm�Hk��0��hvo�q� �KT0u-/2��3�=�2� އ�O �f�])��F[8������X�R7��&(�s�%�R-}���]�i�Tz���*sH��[��x�92"T�GGCb��_��wd��H�P���X�B��`a� ]�LG�7x��ق+�(j��_ ��-����=��mo������A�T��a)_L˶S���e�0�0"���=섒{�P�"�z��ζ]�&�CJ#a����0����!F�<���-W.��i�x�\���6�i[%g�^�γ���t�]le��4GL�?��޺M�f���+-Ԙ��k����$�Q�WT�B@3���$��$�n�u�|lϊ����75 .8i�~k5�Kۈ���8��&�v3����3"��A�x�>�>�J���s�'9��­=������H#�O�a�j'4��9b�����!n��a��d��.��n'� ��6�9�Y|QC�p>GK����[�/���P,�- �M���������}c<��[�	9���7�ӆ}~�r�]fr��¹},r�K���'nP�0R�%���^��;O���fe�U�5��m��Z�~g�O�� �.�ZbN�Y�$�"�8P�f�Mt���-�������NƳYv�83|�U�L���iο�Áo�j6�q,r��0*�Eo��","r��M���	�X�ؿ�'
> �Qs�+�`&�F���D�R$'}�����+EZ�޲�c�._0]Ϲ_/wvJ:ۈ0�ަXn���V	F�ŒO^9;ٌ9�$P�@!Y_B�����IX�g�2��v�b+z3L��u��d{�u��.^�C �7qC��7���{c� ��Ń�X��x�l���d���5��B�|����B2H�,<n_��E�����S���Q`B�!�]}�S佌�ow-�Z�ø(�d��t$6��V�5����0��nB0�(��%鹷��S������/+�^�/TG�}���`Lf�6o7�Nr���$~L@y	��@�Zԇ��RS�񁭧w�rI8���������)�p��t����?F�@ZE~�BƑ����YW$�� ��1�n�D~#�x������ȑ��L�e'J��߉�s�F� ���ǭ;9�G�q���_w1�4Y�-�d�$~%l��n��~�R��N�#`}?���S��4H<��T��AS1���n�WaҎ�5=�k]������MW���+���C��cg֍@`eH��M /�R�@��W���f�heqz�$��˙��m

 _D}E�x����O5؜!)k�B���b�P�Pth|�b0��N��� �K���n���1!^��I���g�&̹��~���.��E��!Ǭ��M�d[b<�����֢���=���般�c�<��R�����0V�_)�:��f��_1d�Av#ГW̘�j�Z���=������,k�(�������2����a��0��cB��V
2n=zCy����Q�'0����{�g���%'K�����:��Cj��i���N���������OG�����q�r;�C�UA�"$[Q��~��1� ��/�O��nu�ؖ]�$(���Kbf�`�۲$��&����*��01Z�B2��3�vZ��o���U�iP	�����i���Hm"�*�Hr�O�z�������b��8x��(�^4��89f⩉�6]؏:�5�(�{G��p��>e�>��p�7��@�L��m�O*S1���N�\��(F�����������B�^+�fo��;M�̎�P�K�̱�gW6Э���Og���