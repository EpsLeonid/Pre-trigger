XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"=�|$���UNlw����P���!X�������b��y�D6���iT��{.�,h�j�5�m����L���5��9�CY vZ����EEu��XA��&�w�W)��>����G�3N�6�]���e�̡˧�Q��`i��r7x.#��& ��x[f��6Ɯ�x>�)_�,q������f( �mPߪ���&Ka�*���k��t� |'.2Jj�����V��b�+v}��8'�`�����{դ�;y�gl-�SYe���Q�i�`���>�Gn7~���eK��f�89yVۘ{n��#�~�w�3�R{%g���4���L�D5'h�D������-'��#�����  #h͐}��sT�^����z�Ƚ�\�*p�i�
X�g�W�s*
4��Q�����y�
k�����p�mѓ7V�l�4�Y�W�?�'%yٮm�w4:"��F�ݜe�g(�����W�������PI��Sb3YE�QR��vl؇��WA �#)
�����˙��W�8���& ��/֫�ٲ��gd/(>��,=�F��5ae�Z��q`�io�#���A����RQ5�Sm��D��'	��e�d�M�����;��(cF{����  ��	~f^𫁄���.R�L|]=u��ݦ7H)ENʧ�}ɻ΄!iEK8^��b���25��6�)+�Ѯ�#%?X���l���S}h��������GJ0,$4�j8���A3�C/=5&��$���&�z
h�yXlxVHYEB    6ff5    1760�T/S�U��%y�eǤ=,?��?���E�O݅{�ڽ�iȂ��R){xo��ʋO�\0��&{��c`����S��q�UL��<�dv�Hy0^;��"T�ǐB�}����Q��?�3���m��=G>0Y1F�(F?
Ք����Q7�l�K�@�{�5s�!(,r%���>=H~�O��ȃi`HG�O6Fv� $�t�j�e�9�.ê���Dy���2�8	�rVBO���0~��_9���*�1��F�������(�w;�O�Q�O,�KVK5ғ�z���T��gB��i�Y�z���>����, ����u�t���E	v�DݙE��@�ك<��7���3e�1����Q�[�Tj��0!�gK�<�u��:M��%�$�Mx��i1g;׮��f�ۛ'_��]A,[9�~#�������ǼMѷ�7��dbj-�Jп���<F*�����=��@R(a�
291T���k.,���φ5r.S����,<��{_}�"�]d�'�%�`����k���[7�e����MQw�^�13���eR=Tjx�=\S��Jù�;��Dvs�*��e=�zǌF����Mvq �H�h��w|�^�eVA<k��3E0j�E���ݓ�CM��	Ѽj}�'�^��� ܵ�8h�!�P�@��
�KO+�M6�z<e
҇F�̽�A��6��� �*I����s�o3Tb$�i�:�
�7����Agz�h�8J"y{s#�!Lu�f�>����:���Z��g��!����+
^����/�ݢ��M#Jj~�)h����i���~�ߧ�-�sL��`��㠭���m@�j:P�}=��K7>S)A0%���b	�7(ʡH��D2��'n�ѢgZ}�g��_�d9��$����`�����CY&�#�b����!{<r�L���9KUSL������`ÙɅpk$�:f=�^��XBϋ"1��MK�+9�=�p�	�=%/,e�_����Ab1I��I"�#4�PĂ�\*H�b,:x=��p�`{�H�3]x����=������oj�i��9�P1��ீ�B�DMNgZy��/;E���N�!����3-� �#x	��r�C�F�e!?k˜%���2O���G|���!�.��0.WC��n����ƾbR���d�W�k[�</	 ͇Dئ3EN[���vL2�N�j[K%�0`=�'��-d"��	:� �P�"c��nu5����'G���؋	3S��m�*�f��+Z�Jp0Z�B,ng��VCˍ��F!��(טr��0F�f�����l̎O�^r�]C��0�@�ӵ���D*:���ߔ��-X��Q�AR��*z���r��cfM�ݝ�LrD�@�G�N�ޣ�]D�ˍy4�㷣�i�]?�N�(Cdn2�l�Y �iZRP�1^>�uX�*�����]�Рd�������F\��=�3\b�%�\�i��0�6���j �IvHAh��0 �dh��1>e��z�1׏��&&&Bi)mDO`�nqD<0B~�����{����B�,P:�S��t&�ʛ��I��Bf�)�������i�%��7���z�!��5���.E3��"s��y+T�&�(�o��mھJ������y��5l�<�#��>(h/�I��幧�Q��d���{���:AR*ʠ#H��y%"|l�^�tT׵���ɾ=���W��B��\zn������ߗ�-���+����X���t�U��J�
~F_cᓟ?M�Eg?��KL�����?PO;S���7��K{�dijkw�!t8��U�T�,���h2��o�?$�8�����Ck�px���N�.��+C�E��Ԗ|��� \ό���yz��u��X�DC�������HS`G����� ���;w,���e0uAfX�:��"�L�J��G�{o�<y����o�X�5�y�EF��F����a�F)��vE��?�'�E���U��B.hW����5SP�u �h��v����߷���� ���b���BuM���}0�/�!!("W�����De�V��K�s���FF��QE$�e!R��f���~C�S�4��-ql]���&6|@K�U|��2!Y�C��b��ȼ(�y�[2
|�p�w���uN����s��5�[b��,�öuR1��n_^��>	���ʇ��K4(�|�G�|O�زfƟl�vN�o��l��{��`v�Fu{���q7e�eӵA�_9���4��|�+��O����$��M-.�('����%�=�d��2���=�,���.�����_�ng�w%�[�TH=��.��%�[z��h��s��X�,hs�<>���#
������ң���F�1t��i� :d�^�]�)M�^m���j�1���A�e9��'����8�)�B���t��$=D�U$�u��?��	D�c�.�2�c����T��X��	 �늻^K*3�������y��t d@.)�a���pO��e����;�l�!������v�Ȼ ��L��wg! B����K�ÏL/�q�c!3��v����s��[�t�~�(�
ۘmg�˩>ħ����*]i#�`��^	(S���W6�4G�<֝� �����FH���bun]��Hdʻͅ7р�=u��h�{�O� ���B��7e�?N(�"#�הr,�L�KͨD;H^�=M��̗�!��f�m�'�����Ȏ���H0/$	��2�q�Oc�H��;���Z;�V�L�6����r��X���禃�cV܈ M�+MMOP+!#(WD�8�O�#������ �(/G�>.Y�P�K����T������&�Mc%�k�mD���ȃ0�>�:����Jf<�F�Ǣ�ea�����>&v�[w|C-U�Խ� ��U(�օ�hR17�1X�f�[�C1���n4�yy6�fF~b�s}0�����7$�ֲ�EvzFd�hs
�DF�
 :k��Aq�|���P{fD�
؃?F1oc���Ed����(���T�\�}|x�L��I�
e�����
~�
4,�>/v��8W!�Bg���dL	��a�g���Ѐ9� Q0j��]W�I�d���?x��J���])�"�qs�u��YV��o�vu�r[��uQ�O2QLo(+�IP@\��?W�+�'��T�F�|��&���Y|��d ���w�f?�p2 }����@�Ӽ�
��JMC��0�,z�6�y��^������N�(8k�
��^%2M߳��Ԗ�{W�o9F��m�ݸ��.�J��5�������>bD���(��b��w�ɚr�gfi��"hWP���N�t�46_�PFq3���>;6�B(�ȵ��V�c�Z�~=�Wu����	���q�]etw�����{�Sk3��}�^4R�m����k^��b=N��#d�'2�EO!E�n�<G�����Dh��A�H�f�#S�K�h?āh�y�~�5)��Ղ�G��	T�7���������rn��"&L䡸��8|nw�|Na�i�m�r�����$���w{�(��8��k�st"+�����J��y�u�I�������}����>?W�c1*�T3N �ȷ�<��b�/����*C"=��(�����Nh���=y��%�$�����z�!��J�ms�c��[dI"�|m���7;�ƪ�� G�M�k�Y��+f�>b���({DH��>�������!(��ܵ|3ĉi�������e�>t���ங�,k.�K#/B?3��|��?��)+\x��|�?�D#]�z7ƚt��6�s3�&z"!�J1
3�L.���d�����{��ۗ	pB�p�����@�����y!�	\�n8W�P	�A���Li�R����)hі;���2y�?g"�&3�9(꡾��u����o�<˼4�t�	�޿b�H )9�6�zD��_L٘�a��e�#�Kab�T�.�C	;$�ӏ�w������=�O��0����7�����w�V��&*�܇���ג[+&@�k��ė���w&��Gj�kg]�:e��@�氙O���SyF�0{H���X�p������"�����eȶ�S����Z=��@�-����q���Ϛ߼W����Ɖt��Y��|��|��j%s�bNzV'����$o����ѣ��J��<iO� \w-�\!��C����'��wtXCF\������>����r4�A�	����`�}$EA=��6=����y+P�N�b��1�ӑ�T�rc'W]�T�p����7�^ڜ^I��G��q!"��E�[#u�"��������}���V��c���z�di8B�.ܣ�Q�ڬ1J����MR�њ�]5�@w�2��$�x_�+�-���8�w���	_L�!�G��,6�ݓTl���M��}�`ɹ0���S.�VFvX�ӻ'Y#������B���*��k/�ozT��Cү6iə���6Hy(��X�Tĭ|�o^����q�2TC����^�����3�r_�g�p�0@N����6��M���^RU��ȳTB�"�{-�)�:Z�M��w����/wCk�I�LV�%ј��7���,���c��!�P�+eNaʝR`�����վ$����r��5W�
�Cb
'��[�5%��D(����v'_"G*�7�n= 8�A�;��"2�ǐ��Tb����n�)VQK��E���k���U3f*�{؎�-9�Vbl�.�<���ʇ�`3�`�<6�Z9��-3����E�MQ��/�n��+bUo�����!��7�ȧ#3����T�&���a��b�rg5�a��S����Ă�����{qY�Ҿ�͊g?Kz$����f9��'��|M��0��jQ�����h��Ͱ���ǒ��֧���؀�����_G�����8�����W/IƩ0I/�'^v�6ʳH
AhPե΄�}>>�<.�����j0�j��6a>�i�)����a~���}�U��&�U����s����5N��1��=B�Q	oTq���UPynt�a��%[z��j����i�����Z�S�tw�|��>���dD���ˏ��,�S���q���VC���c���gJ�D��K���6BC� 0�j><�(���ˆ�u$����U{�+u9R��*��.�/
*�_j~"W<�l��%�A�+���x68�[���g+�k�,є��U�܎!h�h{^��X�}4�0
����lv#$�$���G��~��dC�\xD$6�_���n�R� 2tկ>���C�����P��2�E�κ��Dn��>�(;��<H6�\τ�Z�6�"�d�	S�2b�:_� ���ұ�S;�I�@���<K"���f�i;nغ�̫޾ u��*C�{U�!�RUa���l�Z$�B�"�8��x>��w�������+���H�t<Gv@d,T4�g%ஶ;�߽&��2�'.d	�V�8m�9�R���a6�Ѭ��Ȭ��7m�&B��]�G���=9��#�`f�\�b!�����I	p�{��?G�H3 \��_Y�#J��g��,�)ص��(8qx;s�>�����&1��Ֆ�^��R���~=��d�;��J��sʠ���n*h
Ŀm�r�i�����sB��~�8��mWZ�;�o�(bomw�yA�����2/�ر��Q	Lc	<�5��Nz��h�$��B7�|X}��+����Qx(����jH��s$�A}xSVg�̶ΉL��@^c\��Sյ���Zbc�aא7c �'7�_%#���Y��w86߈i֭�}!�F�u�k�d�U/��
 ��}��cN�Ɵ�I��;�SZ�k�d��Z��a�J��R���?!<F�ˋQD��^�t��������˘>������9xBQ�?B�@���y-l,������Dt��Չ�&K�T�佚>(AV���