XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���5D�;W�*jV���Sg$��2���'pX�y���Kb6�3d��#V�+gHN ����*��.�ˉ|��ڌa�'�]���-m�vƷ��{[�:@��Y7n9��(���d���(N��kE`�0TJ͐���:@Y�+�����;gG��r5�g1+�a[�̚��ޱ���p��VF#6��^=�恴��!���%Zd}=��:'|���d���`��H[�r�W�Ae�ab����:�Y-��{�s��7���'�[	�zE���
"'}�ls�VI���zL&�Z�󯽩�TgZ�Y��h�	���n;���Y���ړCE�����t��7[��q�*x�[�0m��r���-E��Pd1B���1	Byo����/���<Q�a[^�f�$/�J
���j��J
4��p�t,��,y�X=It`��]�o^H9�X��g;�6tA�W�����<�O�VMs�ˁ� sܯ9��2Z7�ل��yu�݄w+]�����y�]㘮����id��#^���-�`<���"!�9�m���d��jɌu������"�vpx�gt�9>ezDx"�GG6�4WEp��/�>G��?G���V�M#G��_#zBK���[�9͸Ԅ"CS��mjHN�-��ɰU���~� O�;h�(uv�˃�4G�d",�{�Nx43��Ug�l�#i:#i$2���%�2U$^�^��<���^�~x_� J6�jy_֡D��DR��h�G�K{J���T^gĖ�yz��O��ɥ6XlxVHYEB    1854     8a0ei��-���^^~��7(�����T3˼�7�lg�VVM凕���C�L9n�"��\7�F�/�|��N���{����� /�����Z��I	���!Ӏ�s�B�n'��97�L�m��sN���AHN�!�3̴��y?].[#�����Q����X[��xƴ1�+���5$���}�-���􇓓�G_�6�2ߦ���B��J+�n�]�'��ت��U:�Z�'�h���?��A��]�D0&�ű�W��@.���k��3s�3H2m^ԡ�_��?����	���#'U)Ch2m���&�0>�ŐB�;?b��]���|J�7�v6�${j��I�I��
jrW�c��y�-ЋiZ����Ͳն�d3��� da���7��u����-SO��#�Ph%��ְn԰��ȮON�� "�!n E~��QL@���=C�e��N`��6���K�9�u�c2M>.��i�?�w��A�:����o�V6���7��0x}��\MVgf��b�l(/a��f�it�$t�i�oF&2&�>��d�Y�^�)���_����t���D�o�rjb��-��ٛ#���Ƿ�����b�f��/�4�>	/`�n<(_��G<*J�����J�jy����B� �k��'c�m���y'��1g����zBpb�u�ټ��ʝ��f�g���<�O�x�.�p�H:�c��N�����+#E��DCK+{�Rʏ���OMW�gf51��9.s`��J�����y/����D�S�u;&�>��n�|�/#f4���{A"/9A�/���W���ө���c?<4�0���q���>/`�4/GQ��T�EB��j�f4u� ύ����a�vSsV��2M}+m�\$4�o�t�x1��̮
1��uXPo�I�6Ҥ� i[���΁'@�Jp!f[4����O��,�T�����9$�PG��ˋ�.]4��ÕǠ�	]?ܓ��uT	���~U&C����	7�y��rQ���/{g��%z�ꃀSf�ލʝ؍�k��?'�$}��7�F�t_w܍K�P�{� 	��|��c)����$�ȫ�;O6��}�I�iFl_+t�Pv�Ì��w	�ԸbB;�J��ܯǦ���b$40�J,r�n����f���������P(ڼ��.��n'��D������"���{�X�:���3����{�z:r1���ETAѓ�mq�%M#�4UL���0:n87Vp��_���Y�ظ�@��q�����M��Qs������y
~oH}�둶�},@�b�&q�5�7�p��ع�-�CUPf%�S�|����
T(�0.|Ʒ��.�;M,?N'x�7�7�&v>�߷� ����ϭ?�@�nػq��L�FZ={��dsO���1�ӯ�U@A�g��9�R�<U}T�����7f�M_�z3*�Ke�{\R���iQ������<�ޠ���-�`Aa��b�Qcޒ����W����9�?�!ų��A�I�V5y�?!XŻX:�� ��0�cs����A������ ������qe����P���ś
�o6� Vz�*aI�a���T}7�Wu],�H�"z=�h֗�Y�=�5[��]`�����39����«�حlm��d�YXգ����`��^#�Yx"�����C�G�U�ɘp	�alՒ��	6��@�,����]��?�rY��_�;l��te���&7J{�}]þ�m�A0�߲�Q�o싦�&H��R�Gv_-�(ڶA"Y�N�r*�+�}���ax1����<n��0��'�DwA������v�e]�;kk���7�W!c[(Cl��A����y���m�D���
LS'���lY=Z���bN�c��)9�J,�@��������u��<�����mPخ=(D*�c������A�:�v06�D��zÀ�w�18}8q8�YY��we��E-2A�ٽ��6�h��)6s�.n:��0#8=J�a��68?ipZ�+��i�hAl�TrCf�঩���,�-�Jɧ� �-�Zbf����e��F��є2�l?W�`>���Z����1���x@kc�u�p�s���#�\C58���t��u��!$��W2%����lϼ�,z]L�F�9 Yqu��`���61��1�~ �h�.�n��y;������/��d(�%}.��qI�:�F��?��QE