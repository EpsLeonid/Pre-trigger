XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H/����mk��{}9;�K� �8m@�i�w�N��ol:���H�I"x|hA��*�npGS��7A��D
ɾ���5e���@��hf#�cPfr	��Φr�N�G��-�9	Ȑ��+�Ԙ]�G�:VD���V���5�@�Y�������Nѯ�%z�7VE�*�����*���s%v��.�^�m%�®�0ٖ=;	�D~;n�i�H� ���X��9'��g{#�<�gc�
L���j �����I!o.�a��l�P�3�I&[��C^@L�������hR'�"K����ɢL�	�!�ob�j~_m��#=�
��FJ{�1�!'Kx���xˢ�5Xh�[�ް���K��0�M�%'���2�'d/�,�&j[��ـ2b�X���٤�MAWm+Hw�	�J�D��x����}	�y�$/��Z҅{�D	��f��3�h�y�w&w)�
�,�}��
�8�����x�������P������s�,�q.�d��W�
� ]�\�:�� ����N��4�5ƀ��ٹWl��_;����d�fL���)��"&R���D�����*Q�" ���'}�h��a�q#Mo�?�~�r%W��Qڮ�Qi���nkO�v���:�%�ϓ&�USÿ��nyee
SQ�i߽HϬ(��j��jD ÿ�g��2�ѹ�r��*� ��Z���!|��],�s�4E�+�Xk#����<��˦=S�B��� 6[z�P��%b�jb������D�sY�%���c���!�HXlxVHYEB    bc57    27e0r%��$B^@'bA�w}�08l��I%P8LFՇ:��2�������t�@���R�|Sb5�Sd@��S���Ae��/}yw���d��-�SS��q����E��G�T��L�u�1�,�O��E��n�V׽c��1��bg�*�/�ʌ�Š`��i�xm}G_(A������3�k4�����d�jC���'!��$y�ןe\W�9�����7�ۏ�vP4|K{9���=�vF��44~�M��>��'H�{~�N�����ª,���o��*8�TJ�	��u�R�uA��iw�j#~t�
�B|e~�U&�!��g0��@[ ����#[���+a����V��S�~Η�$�L0��C�b��T-��#L5"�	��Tޒ4}��!�z�з/3%���NMʂ���,&��x�
�H*˒7�_���CD����#�[~M��z��Y����;Y�6Gb^��[~3��-Ұ�A���ųq���a(�6i�z��9�W����1�q�
�<���1���խ>G�)��d3�#���2Ͱ$i3��ϭWdB�u����.�oJ�b�\	̆9��Ґ�	-X�\:�3��:�����b��D�+�1F�u��_	����KF�g�bǥ�ly�,���A_�t&�=���(��u�H��)��|��1��n��irj>AX[�i�@6c�fI]3H%g�B	��Ҝ�܁$ע��Ą3.�4ߣ54��#���8Y��Z��+Y��n'��A��rp�_j�p���'����t'�_A��τx^�|�9HY���*�������i
x%�>��+��ȍ�;��¬���B��ǣ�&��/�π�̮u����Y$�w!j�I��;�E�8���M<�<����bڙ]�9cb[,/F�մї`�H�н��n�!
�˼���c>�Y���0�f������閼�#>R���d�|6`4���I�g�T;b%!�Q�z��/���>ϋ�V�GO�\Mu[|I*k��أD)�~r��p��[O�U/�����:F?x��S.)��.�N�7���x�- ����}l]m���Q���BGj�l,��ׂZ2N�i��PQm^��:���C�������8��@��0/���.�y!�n4���2!�C��y�ҖD�m���]�?"�C���A���5|j���X:3:�����ΎԷ�0��M�/�4��,���IW@�^�  |�A*�ߏa�ӎ�S�,��h��;\�F�GI�`5��<2֭s��Zr�It�S�ߞ�ls�)�3�����^���C�m���	��[����:��~����4'�R��|��v�"lj5����g����x�\~t�u��Z���	\eFe|������Y�<Hzh�]�%��0O[�����XL4�@	��-��CY��U�l���4'�g��9%����'E�T!�ɏ>����uy(t�����U�[�?;3:b�Zg�"Q@�z�vД93 ���>�ZaMPuݚ�����1�t��f/�ȫ.�U�8��To���~�ٟ0b�#X���sl�7. o�k5�̟$�[��a �]J|�7k�7~�;R�4�eF�hω�R�yA&<���i���i��wcR�RL2�kG��R1�іY��M��4�O$�f�Xε���u�%�'�̆K�������ڍ������"o���ڐ�#:P��KV���=�"k�\���SV��DD7� �β�|W���׸4�AU�m�C~9�I�y�xtO�?�Y����?�:ۛ�)nw8G��	��,U`�����;�
B�]Dʅ1��O��c˱֖��������J(]D|���Ow��7�hq��W pP�Z˨����x	I�2�yu���NX��ĉ���f�@��_2�"<O3��Y�3v�/ {0��$�1�W3��"P�� �� ��5�֓X-���g���jX]��of���� Ay��}$%���q�v��1��I�ks�;$V?J�p�;�&�����}�b�S�)�#<�c�_8��R�4PR�bM���vn����#A����K� �G��D��d��I����Rrv�.�s���β��훸0,�>"�W"K!\�#�
=M�6'��C��\wuGa�(�G�����p�b���.��Ϧ��GwML�2̎�b<܌?LW�$�R�Pv�����^lDh��.%x��Zoy�%g:����*O�S�f8ݤ� D "+Hp�T�r�@yC���o9<\��E������^A���S�������+lu�kNg�,�|ej7�s�!�̦�qج����|�
��L�u��f� i���w�C����(�*��w[��5�wϏ������uh(�HJJ�*/n�	��4#�6��Zk�ڵ=�w|�F�����A��U�F�V/�`�O �ǅ->�G�����Nᥢ �%��;��ۈ�Mןϼ��nP���.��'u� J2Xȼ�sZ#�7�Ba|�6��+cψS��M<�ҙb�7]��>(\D^���K���B1|>ao�m6ԡ˂�⥚�Q�a�&'�\%����_B:���'��6�sʁ��o�Z��7)�o�<7O}{�X�<�pxM|=n��䚴Q��\*uV�:lWl�����0Tr�O<�I��!,�_qCUZ.��8������C�Eu6F���̜��5m8m�*��+�B�H1_t���;�X�Z:M;l)�gS8o1���|N��B�� �{���R�톱��3�n[�
ى0'�!�0<8�ǜ�/����B%�0W��D%�$�2�>�K�w�Ү��>�2��@GP?j_�.� n1ݶ+��H#4�p)��}'�e8�\��_]3	f�.�b,�֩B�t�2#�����Oj�|�CoQ�UmU�d��-q(��[&�A����t�.)+M����M�� `�+el���r{~<���:'}K<e=�]Z��7鿃�)�];��pN>ڞ,�}}���K",���8W;���������T������Pj�$ףx��!�����^|���b(�`ro��$�GF���6s����C��L݄��t߳K�2�[s����7���H�ア�_l��9]��}�!N��|2F��7A�͋����� �˘h!J	Fb=Z��<��U!E��>|č��O�A<�C�s�_)Z�⥲Mt��VzV�'�9!�k#bXn����j��;���U4f�����4�fǙy�pd '9��B�b��Z|G�N�M���������Ko����:�.�i1Ͳ�lP���>�a�;p焧�1\|R��E��Qa�E��WFFg�j:Ig$��=G6b�e�r1�#gopKk�I7GML�K:�u�,Ek�5�Q:�0��Gǈ����A��$$���4�к&��V��N-�"c$0e2�֔0�����4����
{��3z�"ދU�>���<�H��1��ZM0,�Ms3OJ�@�!'L���C-l��Y0�/&"|����%�z�VT�2��h��w�t���д�T���b��X2�k�l����=�fU~�h%��DZ�$�{"E+n����� ��dy�{c2�,��y�z���B�TM&�������a�Z��nٻ�����Dh��Cٱz$ܓ'�iη�~"m ��Tf��������b��������El�W�d��2�L=Fi������jr6%�����]fKMZ���FU��}?�Ud��'H��	>%4[S�OD��� j����@�iRVњUƞپ5nU��A`��-8>���YA�I����HH=+����榏�J���L��-���&�"�[�Ó�aæ~6~��Zd0O��d�˝9U�ǁv��#^�1W��'�.�c�et[��z�t�_�=��F?',n��T�d0&��8���,�\@��rg��q_{��j{�h�6�[���H��%�E��ce2&�6�t2��3�����:�����tQ�C����3lt<^�Jr��Yj)�c �����	���|z?�r⎀�Q����6hѩ��z@y�*8^U
SFX�^v�@�2b Xc�H��,7Jۅ�N �~|=�c����ؑn�=9"�(<�"xbn�����Lnq,�����=c���qB�(�N(l�����&.��۾:$��h�]������͵W%�b��%h��I{>kJY��\i�݆��{�4�L~C�*�=s�%�` =��� x��|%֥{@�T�q;�0^.}�ZAىdR*�n]���
�V�i5Ȃ�t����`OT�����]V�v���@|!&���׍��_?�.�����2�����-�=ώ�V�d���S�j�P�W���Km,�kL��&�)�r_�k�v"�U�f.46#��jU�Ӏ�;q�>0!�ր�X�P�>xz](�D�."��m3p:f�j!w'8�p /-�R����j=T�ᯃ�bD�{f�e("t���1)�J�t���Gu�qW? �-��䈎H"S���#���6�����jAA�)E��/!@[]�#f��*�TYA~9!�iܨ|��Gi$y�dY�BIP�c����3�M�q��(d���6��JCC9t3���hd���X�cp�i��x,B.F'�`���B��J�{��8Q�g�@�j��]�zt�&oC������$�c]�%�*�i�%�)�+�{�t����޼��Y�Ƴ�)J̩��^LD����b�����b���bZ��!O�7�Dnr�\WϦ㯊^���d�jmc�|l��Yb�Lvѣe"6���=��+�ŏil�Qe��S������]�YK�zZ�XޯW*MڂAkx)�;�oU2oj��L=3\��Ao��q�bc��o�i�>��2�p��eg���~����%co	��ȩ	��M1��H�Nn]�?���$���ޛ��2�Ў��h��C��d�u�dv3��1VB'�^O��"x��p$��q�%�����͇o��e�je�V-���������_f������+�������l?>���5/�t]�O�a�;@ D��.]�|C���A$�0��Vް��R�ۧ��c�P�����۩SNW�{a�z������S��?�zԹ �⏧��zϊ@���������x	�aM��	�c�qS��3��&݆f�Nܰtm�kqL� �vd�Gg�����)�HX�z�<��L>4�����L}�n���A����Eم�ҹ3g@y{���䱠G�p|5<WXd��v�O��Cz���V�y�r�`�a��a���v���z~o�a�Q��3��� ��iez�%��a������5� �%:@�+����N~E�\r�W6w+������N� �8lK�#U��ՙJ$) �����x��vP�!�h�9�:^�	�d'�f�t&�C�����M��<oy�_�a:nAm�x ���הG�:�1�!y=?�XV.c5G���	fQ�-^tR��\6w�@�ձ ��q���'��
�����si�6�`T��}�v]+�1-|T� ��E�c8�:՟s~*\�H���Q�2#���!lZ���5<|��9�LZ�mY�{�^�3T�QWu���������q�ެ���fa��F��#��r�Q�v��_[d��S������PB���PJ�>��V����`_���DJ���Q�Ygr���Nyqg$FS�Z��� jW1���:��{���N�w�gPc@���7�MJCAap��$����fXH��9����5�I�`%�_�}I5*���k��V����g��N����N��Q����[-���4�7bY�޳�Z�4�:8����C	�%E�����@�������4׉s�����e�B��r^F���]�u�ߘ���y����Σ/c=u�*on����UhC�^&B�^RN	˸V>��K����|��C����2�e���%/��̈���خՉ����͕��\��?o	'y	$�/.%������q*:�ς��s�F��~�D$��z1�Xßjr��h '��ׁO��Z�V�i�p���~�Y9�3���g��`J�VQ�̟�mSS0�-���ه-{�9�9�����*��Y����˾e�d�&�*,�1Rލh��Rw��,ݍ�/R��uW��Ft5��̊�R��T1�/� �YE3�A5�ށ>L���Es_�Y�`[�/�"~Ӊb(�ѐ��À~�\���!b���fp2�_9�T�QusZll>LCj �$��^T0/899ӐIU��>X�T���ഗ�l\�D?-��C6�)HH��$й�yeaI�
�&��z�d��[5D)�+����&�-�GP
z
�@�w���|�����@�Ω�Tٰ�
��kI�8���De.����>9NܕS���ַ�W���@/;RY�ƫ�2�KFH�k��y[����ff4_I�}����_���u[��w1)�U�06__`ctԴ��s?�P3�e�8���QZ���҆P��:��u������*slhR��h��+5�2$��%A$�<�}�|,�S�h��ԛ��r�:�&E��]I�=� ;�& �x�(�6�V�" ����Vdt����'�Oo5(��f6 ��7�I���e;k-�8�_.�$������>�q?"�d-�4��녓��FbB��
���ȚS�)7�����9���)���Er�UhP��LN�(|)�G�}4��:^RA��q��#"�C�@\݉9��C�I��I�R˔�4A@���Z�5��d��m����7�0G�R�N�ߑ5n��iJ˟��� �Nq����}7�T�A"Ə �sWգ6m���O��[C0	��6wU��kxI0�l���b& ��l�k�}�A����	�I�K ��UEX��HI����	�7l�n�U+�:�xiG��E�(���w��c{�$a7�4l���"���I���	�8%#l�`W;�$��p���@�; &
��3VxV������*I�h
��9�`Xy���}��D�����6�\TU:�I�K�Lb�����L61J��s�ǔxQ�Q���)ÆwX5ZJ��Q���ڌ��{{8!mP�͑��A'"TV@�g��8&��7+^����pEp���0�6��	�{�н���f�=���B��￻#����f^�nd�^��-}FKmw,���Dݨ^�J�6�Ú܅OU���.GN���RƎhT5��ҭ���h�ȿ��S*%br,q܁D�z�!��qb�*��)�#/;�,F���}:�n�,��O]%n���QU��^/Gs.*����~]Hf�	�O^��?s�o��������J�Qw; �<�{ M��W��4V�\�("�w��rR���k6���Y�&c�}�uE#��j�>d���W얄)�1���B�}���%��'�-���L�|����k-�{���<7ݸ�'_根�m<��R$̇ǌ��[�Ȩ�M�rqAQ�z��� �ˋv�S�a�P����Ơ?�у��Z�<G ߌT@�c�hjڂ~~��)��.�>p��'���9�mS�)F��k���ŋS�#���w���P�e�ƗAͮ��<��'�и]�57w3���ۄ�rj���{l�>/�C�.f���&86��LJ̀;���'c�֧�D�b�1$����g�iG��kfB˧v�R9Xk.��G۹]Z:_"�J�l[K�Py#E�O������� ~cY�\N��Ȟ��"�ƯQiHs���Ay�C ��/��&�˭���3R	�)������ߔ�s�j.������j<�]�
��A�$ǌ�:��g���7נ�%�-��4���b���
5j���Z*����J��o�1maڀ/y�4I"]l�.��hh ױA?�p��3�#��y�-���������V�,��1�.��p�6)��T8~hS�L����F(0���82U3 ��ӑY�>K$m��|�^�ohU*�ÍK�=�"aJtm;�P���i���:�5��v�&���&S�`����F��	�������Z�-�Z���T����l�(=KxN�L��'�|PX����`�Q�v%!���4�ݼ�vj�Ưj�{����g��m@
a��5�L�}�BlJ�ӶJ���r<)C�y�����zj��qL�u�<&Z�Tas��Ͷ#B|���ʿ��,�굛�j�N�[����Ȼ�T��E����6�<�ʽɓ��Y�0�q���-�S��P���7dU�N3\y��>-x��(z�Y�NJ+AY?b݇�ӣ���JQ]'�]�=��w���ˀɺ�"3�'m��͆�����ޏ\��kk��2��f�|�&���2��N�UHZ�ElHMɠ��0�m�4�m:��{4�O��a4T��'oi�a��+�pFx�c��o5��F��<�-�Yb��XwY۾��[�%�ߋ�&�@'X���8�+��?��t�@AZ�KHꎤ�Yݕ7�g�K���q%������/(9T�gK�)?�p�v-Ax'�h����i�'!��I+捝�(lJK��N���f�2ўtk1�
B&emqn����(��묏i)[fWi��54Ɔ3d��K_o��:��!��s�\Z.(������w�T��;׽vo�h��a_��(Gr�����R�J���]/,�=?����NH�V�M����=ٞtߡF���F�P����?/.J`����N���s�>����=�{�Izt"�7!�k�H���d���:>`�԰<S�|����	� �ᗠ����̚k�*�}�fK�	<��I?�į�/<�^B[��+6x�)lVJ�*�C�Kv!���N�+jz�q!aŎ٠��b�M��!+A�	��P���������?�x�7�����ἣn o����L#��f��Ñ���j|�Λ��س��R�qVs�sNLo�� ; �e���0����0�](��7�v�����W��(��/h�������y�5��n���b����91Y,ZOv��I�Ƌa�сXT���3�^�#����e��Ԡr2���d#�D�D@�0�}q[�>cZ��1��M���1G�-T���re��`h4�|���S��{�FҢ2^�sF���j��><]�g���)��A�`�U^0�%L �}2�U������ \��]_���5�:����żX�؈�Mۓa#am?*W{rT�е� χBę`���#�j�Sی�F/����&�����.� a�� �I�L�<5��r���X� ��������{槨R���h�������� ����4J�(m?�Tu���L���v�V�1���io�;t+e�$iv�s�<�jP >&D�?Us��I�Z�Җ[Ӱ@"�$��+���RzI&PHk�u��M��@�~��pq#��8f^��Nu.q=�4E�Y�g��0ztu���W�w���@G��yb�����m2/�52o}cH*2�濃xdf��a"&d�9���ͽS04*|{�U-���@Bg'a����o�=�;`���,��n��<b&ױ�C�� �B��;.�;����͖.ā�U�,I�1V���5�Zt�s[��'��6��W�cɌ�Mz৖�1�>����M�}M��/ f&��3w�����c�d�Z;��9�p߮4�g�D��f:�(L4[�_r�5�i���	���.���*��"S����2�Xh\��ZZ*4�O�A7'e�����J��(�w�����J^^Y�>���n�\{��IoW_<���A)\v ,ĳ����]צ�_�?uW�5t˺i~�\}*Y//�6��:ɭV����H�̺S��X�.�ђ�r���+,IȨ�9���:.�Q-���w^YO�^N�0�A����J�"R�K��u��茷���W�̡�Ne�C~+��5��;@�I?,Ă�i��ʡ��dk�va 3w,�Ĳ�Rv�ȤZ�l�t<�|$r_�u�9�d��B��'^�ꑽ�Z}0�ͪ���΀=�(���4�]��:���H(j�<U��ĩ��wr�ֲ�K�q"��T��=+��gR��N��O��uX1�s��}��\^��������MY�3�%��RR�)��-���C/�U߄���ٕT�gv���0�d