XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����?����N�ƞ*ud���qrj�Tjx��+[��p���l��)�ey��R�k�����|���IQ7����B	t��;�ቋ�Խ�&)�J�j� t+Ģ�$(ovumXg�9�bQ(s��)��ɋ)GQJ�L\���@��*���"��if=�Mq�?oXo���A�$�J]>t�K�+��YpD�����m�A��uVW/��R�9��e�,�?d��l|m$���nθw�j�����|ys �!6{c%>��]Q���\���:GQp�U�E̩��7��	P�W�V�siP�(��pv,��8$�2�Z�m��Փ	~�TC��WG�zG� 	J�<\��C�I��¼��� ����CB��A�����2���؟�|��:A��M_A ��K��0�jy�\λ�2��i����љr��U�E.��"%�l�1T\�B9�)���4��k�m1,����;Gʾ=���!�cjy�U�#-^��TQ�?��Y(����7^�E�*9_f5˗��͞���qF����x�V�D_Vb�0K�ֆ}N)�չ�;���'z*��CT�+P���Ģm��8�2�C�S'��=pP����D<\��G����a����Y�&',u�� ٟ#�3:����4������b�bo��2�/�A2|k��e���{�ě|0�~�v*S���h����l��4EA��ߣ!򍄒:�9|(}�����wc޳�H^;)A5dY�d ^Z�
ڮ^%�HXlxVHYEB    5f5a    1490��¨����9���<�8\��Eb�H�@���*/l��� ��2\��m:�^�ø�}c4P�I��>���Q
��id�y<������h���ECzb8g�jy<������\p�������@C{uTZ �$(@��5�$��\�8ע�@�0 �%0r fn��i����L�2t"xɭ�@v���u�I�1���q^�&����W/�2���s���c�h�|@�L�P %�d�dzS�>��p���Xr������$)=�L,�y�F9#�AX�r¼����h��l4�ncI�U��՞�37
ٳ� ӻ�f�t� 'jjxK���S�gUOtw��Y�z:zq���y �}�c:��%���\�Ѧ+��.�ц�0�쩔MF9�L�׀��E�������%e���f��L��R9�>���d�h	I�+��$q6j}�f��5Zs�lI��L�YK�����"I�����_�v\R/Ĳ=�� ������,�i�%\�0\��G��cLiF`�7T��]���B_%��E.>�=�NpíR�� �{[΃Jl����f��aG���>�Ĵ���^ }8X�%~L�&��$M�:����kT+��){�Ɏjf�:�(�(��u߬հS0�d��Q��aDh��U�Eʣ �|EX��Xxe�o�s�DQ�F���>'-�����D� �m��7��z�,5t���Ot�䅒gq����=ɦ[Z���aa�M`6 ���x��mF���">�'�9���#�kY�۴Ξ!:�d�E����u6+;�vM�>����-�%�e�<4]��;�5�n���|ۓ�^����7W��:n�Zw�f��~]>�ǚ"O��_���XC#y���aV8�W�ma��3��b�/����c�����tp!��%"@WMb�����"M0d�B��7q'S$� �����C���0�g�.� MϣSj��`�ˆ�Z��(JkL��S�l�n�ꁓ�D�RA�c�y%Ǿ��&o�}'�}$��fa�_�OSB��h�R��@�'|�#���d��U� �����s�&�ƕђ2��8���Q=��YΦ�*FIiݖ�������?�;Mo�~�4X]Ckܡ��ڗ'H�A
R�Yɜ�Y�d�h��=��>�'W��_	s��$ּ;L����b&�T�
��*I�Qbk�vP��uC l[x(P��@���?Q}ǥ�U��8(^;]�&K���H�"b�όl*�����־˴��ZB�m�P��;�DY/��9��RA8�Ն^{,�'/{�5�!E,���cq�ᄁ���3�� o�j"�|R�Q�,���CE���:(�r�����?'�M�������K���Y'�d��X.l�YOm���M���~J�	P�1ybO/�{D�S.���d�����aR|f��2��*��;#�C�����ǈo5�1:A��w�J1�{4��ww��?�v&�#9�(MXh+�Er8�,R�GaK!$���"��JMrв�ّWIbt��e�H�ĕ��`��*����i�e������&���Xд>����]�,��g�x#0��ŊN�P���Gq�:��`6�����@���C��aZb���}y:Mae�`Co,, Z��M�ڼ�p I���xb��^sP	)W/�"��M�)��78+����[��jH������Q�,��?pP��p�q�3�G�r]J���hx����B5i��巈4�Gy)���b ��/��TL�@3L��T_���T��ٍ����)��Ȫ��}����	��j��Έu�5��v�/���L��=�����=�t=u��Ѩ��D:*��Ҝ�"Zn���o�Z�s�~��+_�X9I0���� �d"��$�D�@.m�x��P��܄A�����n�ó�r��a���2w4�̬��������q�"IA�-����-]��UT���a���䒄v��)�܈�J�(�WC@��^Ad��]���{{�l�t5�`��C�p�°i�'p(a�� �:�8�zKT���z������&�eB����)�i���,�-����i��q�06���r��J�]���G�LWK�P=t�w�'�n�
��u|��`!Fm8��L+�]e�d��m�����B'��%l�6�k8������8��i��eL�Pm��8t,BL�N��'�I��8��yK�}�E����}C�F��$mѮ.����B���lw.]��TM���Pĝ�fu$���]* �\�!&j�fq���W�!����9��G�}�@:)(�kX�����Fz��?
v�Y�̏p#(b�^AF��̏�D��+��>u	'N�Fd5lꮝ�'�|�a0`{�/�����Vd��蟪Ծ��U�#z�S˩<Z|����0	P������j�c|��<�|<r�}���t쪽��8�<#�U�F"�*��"5��Oܩ��_�ԏ$�o�WsD+o�{aN�a#�2#n���2'�j���3e˰�X#�m(fa��|�g�l�v�f6 �b��4�3�����Q>M�V�NE2y.jj��\����z��?�{�9w^`�_ "��@�/�2>�SR@֤�]��:��&ƞd ��&>� WЅ$���R��)G>@s_"h��]?�N	L9�nD��k��L���k@�2T6]=<G����ɱݼ9�u3���r#^��.��C�긵���m�m��#����	�`[� &�g\�`ɰ-E��a�K��8	.�E��~:qC��(�4�7Yj��T�w�ܦx��OO�Oz�+>�tá������5V�U�Q�pU�<��E0�[��.Z�	^¾�)u�O�������)~���M�M��kή��H�S���c���5�)h�yq`<�{��X�����t�#ɋ��ø���a��:��a�z`nP꧍�߃��]<A�~��ɳ�5���ħ�C��h5�Œ4P#��׍,�K�t�V�H�ע�0Zb1�w_����G��uI(#��q4Y��P�
,�ŻF�p�D]���6������`�)��섇��"�J�ЧtD�g�.���?D�p��A{�Lnb�>���EX�q?H��<
�Ȝ%��E���~����S(�ԩ��\�x�bApާY k����������m� ��J@���.���X��5 e�	К��	�i,ؐ�Y��5�L��8���9��n	��$[�:�-��ߨ�a�x�c����|L-����k_�ɖ6:ׯ�`-H?XL8�����to��Ȯ�Vr$%Ft�H��^)�گ���:��fk(���*2�`�~Mɫ�pO��������Oj7����A�+ُ�����. )���DP��H5�VS8|��0�B���M������$�L�yBO6������i:_x������N�;�N��bg	��� �`�����St28y�qkم	8#�Z�_�迢��3K�A�7g�������{CY·'W����&�h\
�S�¯;��y��\��3��I���*�m�+$Teb�w��G<��5�OG��l���C\8�j�	&��X}8 a�jO���(��	��,f��SS>�p?Q��Ʃ$��D�]
Q1���@j�_�?hx:�QL�ΎWi�q��ݾ��A��8/�7[`�����N�T ��"N�V��K!����c�uI�M�r�Art�O����]>՝�"����S���4"�w2"�l��0���s���n�u�B�RB��]G	v)2��RԮ��<%�|Y��0jrՇ��W{R�X��+�n��6��-6��:bFb��[�=o�zi�F�{H����$�\`���j�~��	���d�踬푠�{�a�(��[�d�Y|�@���;�7�J}������abf��ebÝ@y
YD���5{�&	 �����`'rF��G�z.1�����j3���f�p(K����˷�ᄍT��t��
�����f=�8,�Y�Ӆ�6��q����4�lSCT&"�L}��^a,�y�&)}0E���¯�8?
���W�� ~��x�Z"�1�!{H��o𣹜n�������Ĳi��<���ڧFt���P��t�YQ�A-�1�������� F����TP��뭪(Fb�'=��ISA�7diz���7
^!�l{l1Y�FrԂ3c�F��n ���{�gx��yC:"�Gmܵ)	\g�G�t�h��B���FKC3�Ʀ�T{1 ����%P�r�� �*}�T�m��ј|���_�ȩS�xZ-s��l�b\���I�/�X����p.[��u�>�f9;9塰��-�g>�O����;I��y49:|��U��l06I#�"�d͡ܑ���
QQ��*�M��=O��T�.�y��h�G�h���R0��(�]~�\ !ݏD��%�eK��o��2A3i��8�b2�����rG�Ɓ�����M�j�U�V�;�y�V��x@"�����-u׽Z[���|�rN%�7/LP��r{|(*t �F��[8���T�Ϙ�}<�ȁ�8��p[C8��w8G���ى�BL�ҵ+��kQ���;P�UH@uV4�#��q%�=���[� ��UnC��,�X��GU�ƴ\BlQC9s"�+,U�/qQ�A��YZ7�i���2ʁܞ��2яw`O����VFԚd$�v�����V�� �!��'��%�չ������$t�cjqL 2䜧��nn�u���ִ2��9n��7�6<Ɓ����4�E�Hߑ�m�����'�<	{V��ax��v�W
?Q����2mĻ�&<�L�ېd_�WZ	η�������e�֫G`�w���#�f*��U�u?�5�Z+��Zw����J������0>K�|$���h��7?i��U����~��0�BZ�P�SD"P�xV�8rW2T/��۴��0pzP�x�7�(�!W�89���կ��[�Ƅ��v�X�wz�Ỳ�1n�f��И�/�Z{m�Q���ji~YyQ	���ND}���Τ-������}y�����G�O��/MJz�U6������&G�o��c�A9�� +������ j�ܜ4R�k���֙�TX&�_(�gF�"��7��]»9��_�3�L)\��"z������!P���q��Օ���-/�����HU�[Ro��i4i�0��yg�x�3[o��6<6hb��0��!��$>���,bI�W��^�	̩
��?