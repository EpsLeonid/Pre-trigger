XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|�K.SH�|�Χ���
M�}��\M-���4vʾ)����T���_Ȟ�$��;�_�4�#�9�U����%Ro��q������/H.�����x���o.�8K��"�䐙���b��π�cE��J��y��&����.UD"���(��Hq���e,��N9`Ms�l
<���+G骧ڃT�;d�^/�X������&���洎=6��/����Eڨ2����*�HS�~A\��(�б���z���[|�A�	\�+�)�n�m�D3���d+�{/�%��#\E�2�	��C�p�~Ԕ�i� +�����]��ޢ��*DW��<�GV��]2��\B�����t�g���+�ooKKѢ�6+l�^�N^���*7:<C#N�f�����O��{Zמ�{��+�����l�,��E�X�	8"x�#љ\�~��9�@�"_	>�}��J���i:|�o��!�Ll������j���m��ݱq��MTg�6����=�c����kX�ܢI5I�tm�pa62��ʩE�h}W�����'UDk������8���	����Ї��g�,n���?�;�~�k6w�"O�
�Z�!�����~Ҽ��1H��6� �
]�Dݰ����МFi��E�`M�՝���ա��;"N|Wa.�'v�|L�W�qONzA�'��Rh4Fy�ߧvxX:e�a�p�n��@�$��g�����<�j�* -N�͚���'p��{��f�j'����5�XlxVHYEB    1e12     920�S���]�Bvo�,$y����-��2�=dJ>��;3�z(�B.�nJ�6v�����B�폓B{�TF�i����eC�I\�Y:�B��Y�X��F���X}<� S7���߉ o��.������!k7�UV�*j��t,C*X�*U����Ӹw�q�cGřG[6[����&)]�$��ܤĺ �r;+&p����O��ri�d��ծ"n�ӭES#��)�ۛ􂩛��~��.���]/��S�P�O�q�\�t!d�TD�ᱳm:��1iO�]��O���JY��B��|�"L���6R��0�t�	~?�ah�qTm�B��/c����p���a����C��B��F���z#R4��B>��N���SZd9�?�����VW�kE@��3+:p�������Ǩ�)��ӾR�(��+��֤����}�#�x��˥��dV�a�
	j���O"�u3�mv�Q۳�M�6E����	��DҩX�0`q�Z��~)�y�3�zP��|�Q�\^�����
�4*��I�LgB�s2�1m�s�x���U���;��k�6v���W���z.����Q��;NtNð�2ھ&�<k/�нn����'ȴ�M.�����S�.�E=lX�9� �8��酧w�*-Cz�S��E����a⬬���*�nO\:v��2�HB�m���߾Cƾ�r���rIj��H2�w6���H��TN1��me���۾���,"�x�7�z._�@�Ӆ|�Ձ�X�%!$���bO�L�f�k��y֞>~�=.;����5���k�C�d��=���b<��۳mT8Tf�/�v�Dh�l����^��Ć�����B{���L��[������5��'����)xA�W��3�	���94E�z�L����ߎot�KB;r���.���,rP�F�:�T�G������P��V7;�m�E�L����k'���\��E��ލ8��P�~7�Val��0��f}q����_��h���f}>��+��]����F'#~�/o�<b�hʃ.�[�o�@�c �YS�oL�`@�.���w�;��� ҥ�1R3a[z'�DΜD՜b^��Q`���L�t�	q~@�D��R��)�m�R� �AS`���螲�+/�X~��,�3�m��͚�i����C`<p��oyvlHt&������8T��|rܥFqc`�TV�E2��zp������J�����"�v YG�t���-��\j�<l�Ǒ�Nk�h�W?S!��&=�4f����`�:�c�,�%y�@=�C�1�s���j�i��^vd�<�O@�S�wn�p�>%��:�W׊��C�mg8t�+�N �X����O%�&��+�����oQE�82�Gª����ܜD9�S��9�|5+s�S�\(D��z&4�)|�[&�}�Ώ���Ƅݫ&�J'��9��xlV>ac�7re��)�S)��D�m��r̪�.�zz�Ϟ&Zرc����a-�lQH@�|�2:�:��ޭ�RQҀ���+���Y�a?�m��eƦE��'[�7�V�+W��D8%О빅��<E�g gP$����i�F͘T!4�\����nVf����4n��؂7J��d���|�d�WDo��H+�q���6�I%��o�sj��*�׬@f�tgn�������F�ȫ�����]��4���,���C�?��j��Tl���+s��z4����A��Ξ�Az��p�"��i�7�p�Օ/���_�����i���ƣz�����������`(5P��<���G[�u����G��ώ�I6T�]B���J,`X2�Q��F�<�t]��2�mT �HC�A=�r�QC�����S����5Nh!�х�>�wa�\�04��u� �H�� b����,(�:�
��2FM2�-!U��'��lsޢ��e����rW�D,
h�<�y�Xe8�YrQ�FY�Tn�nK+у�9��f󟫧���e{��mx!�1^�D)s�fVl�d�R�<�g�g�(�=��h��t�H�:N��űv�dZ����)3�l��`Ϡ��] S�>���c��ܭ���p��I3�|��K��ҏ�k%`&Ǫ��~h(?�I�=�6�Z�+�	��F *���������-j���.���|��[Ԡ�̱11޻Q�%%��Ia��q�p`x8E�SAw���!F���������;J0M=�4�HҀ�*�I��W��8T�!z�9�Ig��}��BF�-^*b�K�D��y2F�7mW&(zq�.