XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� ��T�N�!j�����Wa��6c))��:�=Ƙw����i�[������X�����v�ܼ<�{c �Gf�6	\�"QG+��s|���#���Z�j�u�x��lh`}괞���	���%bڝ~<vF�V�k�YÌ\��z"��ss�%C�ݓ���ͽ|��.v��l�2��i�D� �EJ�V��Zy�).��4n��<g>����1}:	@O2~4
��1	d�-������uʩ6r�V;K�����	@�Gt�_�q��̄���,�Y�4 �ȍƙtA�p$�Ͼ�A\������D��ٜwT���! �n&���Z�����1�+�����L�4߮��`�C�g��4��j
���I;!Y�df0��$����Z�����3���7�L8�	6P~p,;��p{F��^t���0x]�ΔKF\�����ȍ�U��ɦ#�^�^*k���y��:˰��S�ԫ@�Y:J���:�D���u'��݋�2#�����삥����hN�W��*��r���-K��3�)Ƃ!41��]8e�7�;��_�uρ/9��j���gɐX1L�aǡjg���19.��+�����F��}l �=�#����	aR}�%f���Ge�B����V�F.����������!�<�t���*�k���/d@����P�ɼ��J��t�
���,�
�l�J>���+�k�uZ��`s������#'�#��?�#Y̋�gW�w0�K����E�F��Y~	,�Qb���^�[6�����XlxVHYEB    fa00    2c50���Z"k%AUFv4�J!�؋��33v}��}^/�A�Svb���q˓��%�+%	����}���cD��f8m<.L���T�R����)F�y� ��m3����e2e�� ���pJ��ж��"W�.V��:削�0�??0�3��*��G�K��_T5�l��?7^	�1�L�ӬH�$s���	i���=K8�X�}�/ �5�i�h+�������� �KQ�����e	Y���.
Uۘo��T6U�dxU�S�w�暼z��\zJ��y�[�ߠ��d���i�Z1�{�����'VD�S^���?FEc���q[������mgtU}G)v�[lqf=��Ѱ坭θ�`�3\$�k�C�,^l!���9<�<=��]�� 
�����b����5��~Y�Ǵ��)�<�?�7��i�O�B�D' x���Z�˰S���46>����Vm>\XrH\��|�eh~���h�F+&~2��(8s�I�y���F�L���{��3p��|��B�l�.v�G�s�d$UǮ,b�c<%
J�I��[!PҞR��>�Fg�q	PW�u[�k�l��_2�
��b������Qm�h�
$J�1�7y{L� ��Ψ�9�[���d�Q�m*Ͽ�7�l)�&�e�a/�] ��d���f76]�[�*�fW\'w#�B6��O�nOX�����KE�Q�X�'G���N������p*w �P�Yy]� E:��#`z�s��t�.���P3�C�\~��z�`z�^�u� ܐ�)A�e��Aa����Z��k>���ˉ�N;��@Z�Ogz ^��Ӷ�ˤ�&�Ͷz��k��o	Z?�D�j�8�}�w�Y��:qy�����6���� 2$�����!�I�ƈ��9+�yE<��c�F�TJ�b��.r��A�g��5��X�O�s�)�X ���5��$��"��-a��������P&�V��%�d2{���Qg;�S_���%@{���?A�4��.m�Qws�CI;}���g��Ai�ju{��pu{t�R!ɱ���H��잢��?PQ���u,$�OSe��j����0���>BK���۷���V ��1�đ<�^�7T��۸b���9&�E�v8#X�ǃ�2e�D��
���&�m�,!����0dcg��0��!tV��e��z/r�
գGq�?jh=u}Ć`���1��τ����UP��-��%h�q�(SE�5�7��0A�tJ��
:�W:��?� �g�L�����\��b��Y*wl��p�AU"�r���]H.*39�1��H�'�F��=y��όn<R���Oy���79��}a���0F�L7϶G�e��S�y�.�'�u��.|��� <�׃2�jo�`ԁ��EE��������9�B$S��0CY�G��W �7�w	�$[~&� %�	�j�@�� !p�=Hg�^��g��������A�����Y�IĖD����G-k|��Z8�a|�C���2-��7ټ^:D)[�L�3h�[Mdc*K�_��H��9�d�6�vx����XE/ql!pN���q��&��a B����������I~P�^�fw��rm���\�G��O}x�N9&�Z����R�P�}�9;j�ۘK=r�2(^�y**)��\�9�Zx ��������5?/�]`H��?�Z��S�Yּi:@�6�(�fB���SU��6�q2#��^ v">�ɗ��8�h�x��n �B螪��w�\�cO���FC %���E���clQ^qC�>����($:��}�I�J�����-�K���FI {�y��2�o�%'�'1s�`�m��#Ɠ����hҀ�� ��ܮ28%�۷�[�b@B1�J����V+��x�������	�L �N<�)��Fʒ��P��Y��A���kˬC�2�4:��k�%��2]���;�Wi����8{GN�>��;�~�N�]z 7c�9�k����&_R_n��B�����,[�j�i�5�7VLȌ��+]�d����K]l�7t�Uv��֖��k�{U\�˙��X��J��45C��:M���Qm�]��������w�m8��SI��U:��u����y�jSJ��F\�5� J��H�7�=�x��%���y���ug��P��n��CBaxR�^DBO�.����u��>6���:g�.��"u���?Bÿ��:I��B�K|EIO���5�NO�h�������_Kt�yRZ��s2� �s���ȕ�"1�2ktda,41g�,�������@w4*�G�G��Jr����D���Ĕ�S�ve��L�Z��_	�\|���1�$�Ky7�u)CD��K����߶J_%��������m2֨'��JO1�4w��C8��ّ�n39��Ɇ�n��k��~[�ҤUv4���i�b��F⢤o����Ҧ>�mi�szȔ}%Q��v����6�>M_Ԟ��2���O������#��O x�[^��#+�v>.ĳ��Lr_�
��N�����q�@Qb�O�R�'�!!�������Q� �vpЦ��`���(�s0�����(�a���F\�ľܵ����ټD���1|S���#4��@�AuO=,��ۢ	N*�x�*���߼RYB�Y{�I&\z�8��}qg�F�s�H��\;G�]�nc�N�#&)b׶���/L�|@��ռ�æ{��|]=�'�0yk�:�|��EQ|�ͯ�Up��n"��r�\;�˓�H���!�@�x�0��K��I��Ӛ���N��2��**�
5t��u�=h5<(N��m��]�xJ<���t�1��F�������cf�r�Z�Ȩ��`�TcfE�O>VZ���3������� ^��yz�'�+>�]tuƁ���n2	��O��S�� H����('ئ�k��EN���\wTY��&�a��71 ���������i�5@�̃H78m3D�fl�Z��F�~_P�Z{r��|���8lX�Z'#=�P:��~�^^��䍻A���F(��Kd����4S�N�-VZ��`��!������`���	y'Z8w�Z�B]q�1o���������݋�|dh�B�F���
��}�9���	=NY[���>9��qIF9��[���Ǹ*�n�q�;u���A��æ�'���ўYM��b�{}�����~up�b���{���FO���|PE��D;p�4B5��5GK��Vɷ��A4/i�YO�4cI�	U��\,��B9�ܨ�&��D�³�������2��kN�i~r�֓>0�ot��YK�F�6�'�+���ݪ#|�������m������G�\�qTմS���RNcXw$���2�$��|P'=޹��=g�6a?\���[kմ�׉@�{'��+4BL�˱�w{<��En0�f�v^��]EW�Ԓ|
 ��2�5��̿`B0^���d˯\�X�`~��o����ՅA�do��ܗDK"�\$pA�H���.3��Rۇ��a
�٫$�5ֻ^ڂ��s^)�[��N/q��hT��x��U�@D?0�8	m��BΟ�&�]9�+�M*�d������M�����W���ı"|�Qm0,}$ˢsoz*8��.�U��.���!��rcS,�%��<�If��V]�� |�_��Ջ���]�0�y�̶��9�f��(^+��K���?	��d�&�4�$ɸ��M#��YiƊ�2aB��F�n���Ǹ^3{q�@`К�C�U*�A�1�/V#������l�4�/��n�t��	Tr�Uh/�p��n��p �������.��A���7��4��\���`����N�PO�ܸ�ͬnk��c1�5�>����ʗ�)�*�HJ;8���W�cq,D�X��Ӏu��P�:���y4���k�n�>�[;.:&�R|�fΏ�<�TM֦���!�I.z��#{h�b�g�N�?�ވ�����m,�y�E��ǚ��#+|�IG��W�g�w�ĉ_�fv4�Q�as8"�;����^�3�C�q4��¨Mn����>4��_ ��Dd��w�x3|�~�Q��ܑ�����j|��+��,]���g
�z^����b���`M8���5[�5')p4���u�	L�7J�rq��bt�2�\�s+o`VHAq�XCV�El`��>�4�X�R�V��ǳcI:��ex�0m�|u�o�.[�%��򊎓Q�(�3���b"+{܉��s��̞z_��{bp��\�n}�	��RĚ��]k��7Νk�3�B r������0F�סWt�|+���6K�F��p�q���O��̫ SjF#IO�tq���t2�^��6BZ��P= �"M�D��9�"��r�fP��s���BذJ���Ǟ:v��i�iF�[��t�s4Q�� ��]�+�N���@�x#�����pu���hx�e������D�j� �w��Q�M����y}95b,��H晄�3E��\�L�4�X�������Pț�3��4�D��[⃑�~�B�_:Tn�}�MC��b��n#�)=Nh%��=����Բ}PH��R-�d��b���/���H��Ө�}Ԡ�TĠv�76�U�c�'��[@�0��+�#>��6���������o�x�!(�φk蒹|4k��>h�l^g��4T����4�}��*	�a%���;�9s��V��u�_2��͵Ǆ?"]5f��10�{�"�/�G� ��8x���-G��xshH/<tw�k����T�z��9A�,U�+�e�'����dܶ�>�ӈ0Z�H���4E_�a���y3��S(1�/��j�mYKj��"	�xX���}x�������<,p�Uf�٧�W�½j��3�b�t@�^��h%ʻtC���CZ1`98F��PN�FS��Mv&��\�Ϡ]�H5��q�j.ԟ���h��� +x}9��p��[�<I�Xix�����!T�����6�%����,���-�u����@��ΚT!�x�����_�1�J��9���_c��|�	��s�����O�=�D����Q�n*q�dJ�e�y���ff�>T��l	�E/��' �@����l9�]8/��)�9��W4Ɛ#�Y�6}�Ye\���ȕ_ț�%S�`.V7W�8��Z��H`�����Pj�4�S���p���㌀HM��rh�!A����<���ӊ��_��
\j-Vġ'�?��C�l�9=��&�E�Bd�W�H���pj8��G�}
뵋��h���2�	Rm�2�����L��kn�Ym{4�03>� Xby�l��C�h���{�, "�!Iŏ�l=�R����)a^)�HS�c'sց��\�Ĝ�U��0Cnl\ 9�ola
���BN* �l�+�����g_P�<��l���ΆN�+xXh;"+ߛRhu;����	�\x�{,j�ܿ��I����F�<<��iil���/��bӹ�? '��SB��RS+�?e��e��������y�JZ�n*=7;{@ؔC˿q��T�I�$>�o$�d��(8�B��`�f��C&�����^�*f�u��3�/����;��u�iNQ�D�<r,�nG��obQר��n�mZ��z�&hi�����M*Q�������=��>L�<�E��N�{t/d�ɜGͲ��_h:����_g�)iK�>[���%��-h�Lgr���4��Mg�rm�����/~����i��6q�<�����0�Y *VN��ܝT�|�������lO��>O��%Y�C��Y=c�w8Ly�A���ZbM&� ��ןJ�D��<�h=�G��֍W��/�N:.��5�2=�_�t�z��RI]��:��Fs~�;�՗��V��� @R"ݨj�F���G�)�,G�p� �b�B����p��Z����U1�՚,GO��� ���"1�� 䧵��5�2n�1�T%F{Z�Ou%@�^L�[�����}�GW�A)9I���9X���E��&+���,���D��L�^Vp����De;-n�/la� ư
Վ*�spJ^��H��0]*s���~�H����)��dc�(����5O�:o����U��۰��#��I�@�m��%��/s�4侤����d�E�$7�;]c:7��7�96�\x�Z86���_���Ėxx�(8��"�.�I���<&~ql��4~��H��)�QEG�0��4�d�I��o2�V��e'��1֥���H��_�݃�e���ZʵE��3��@ԙ'57]����fB��U8Ae}��%z����m9~iOŇ�-�3���	�-�Er�L�"�Y��2�/���ą'��x�w,e1h~N �G
 �}��3�Ӎ��r��H�I�Y+
F'��Ӧ�o*L�$1#G&)�llSz��#i�ƲN~.�l��D�TL��Lf��b=f~�����v8`�â%0F���W=>�
����q�5K��p�}�`]R���+)
�2���ii��O��j��<� �ƼZ�
ъm����0d�U__v��Z���X�%�S�GK�Q/V˩�m�;�Xw7Fk]�M1X�Ʒ�l�Y|͞YUL(��p���Y�s�f̗���QW�ȑ×}a�� _�	>��wq����V�������)�����[H���[�1#[�%��/;z���C�p���RPrn��p�9���|�|���;�o�����ܐxZ����@1oyq1�� b}�����'u/�s��s�IX�L��뢓c
|�� ��19C��oG=�~��,��Ӛ��Q���3-�@���׆�|n�P���\�w�F�����_6<x3��~�LH���!9Cy�%�$_W��D,�)�2��ˆ���I���|l�H�6*��p�g��t��d$���iG�0F�HaL��)~s֫��|�D�Dkٙ����Ew�h��ѩ��0�S:��7h�P� ��oǰ,�-V�:�����\�tS�@_��t�1hCW.mc����#����V���۪��WŰ��#�oa�~�!�AH[>�� ��`��o,�l�';Z�%q���bL!�+;m�JH��w�_c�����n�� �Nq�_6�;�nd���55��S���7v����D�{g� ��d�,�I��O#$��|8bY]�9o�W}�_�M��9t��0ι�%�;���Q���g���ihmo��s�!�eq7�z�7d
aW���0΂ ��m�i�dx>�)����G�B��\M����A�ޝc��$��V�l���k��Q�ؔ��EX�Z�U����C	M���8ʥ *����k�I����vN�Q։6E��£�-~xw�(8����_�m,�>�9��O��j��Ũ��n᫁e�5� C����x�Lц�t F�|��4�׬��	=G;^�� W�5��}��CUt<�����Q+d�i�U_�\t�/|TF�BQ�&�xm����k#�Ͼ�$���q�?a�[�����#��+�^=z9�*A��za	��5F��!D��e	�N�Ć����4E~�#�ӆ���=p��3���˒�|�JF㯾?�E�����VJ^� �rCO,�M�:�L��S�"4_[�f��I��Y�F4P[�`�hħ�,\�F���.�EM>�^�AR�X<G�4��� ��Ry#��A���IrN���޿&jԢ��T�����k���ox�R��z�XXwU�V>(�1KO�υ>��&�kN�X���[�|������Q���F�'eD����nGbT���,�"�6�ٝݑ��cnf%��]_KJ��J��Y����:Z���_7�r�_F�v�H!l�:C����X�{W���õq ہCI�a�'-;���d3A^>��B� z^��ϹG���#eBF �5�8Ш
^�w_��{jg�mP���W!�5�]�Z��=�[}�P�g%�v�)�5S��S�4�nqۇ
n���G��/�C׻؜K�_�|�+Q�������Os?�L�����?�ut/����:�6�pg(�叾V$Ͱ	X��`�ܣA��/ܑ�Tvw��T��?� 4X ����s�>�?H�,s�b�����'�
�<�[طY?Vo�e�"�G��T\��[v -�:�Gt/�0�d�f�£��3�}t�����S��P�z�3X�����,�+��#�\$7����LXў�(K�?c�������RL���!2��'�s-��p�%"��3{�A���D�:~0�Z�����C� i>����)�qN�N}ԙ�"5��%�sأ����R`�8�o�b�x����QEPvgH|��ᙰ�F��� ��
BU���/��g���ɼ�C��z��T�>�\>�v<@���'T�k�{L&q����Q�+� ��� ����FӿR��Y2x �S��d)�E`���	T��r�a����ڰ�C�A8-�_Ws��z>�&��|��:�>�;���]�^be!��F�"v�<�_�Q�:�Z�H�8/֋�����qx�"�v�ؓv�[~��� O@~��)�^{�:=�j�-S����,��3���dZ�I�ZUC����v{��YT�p�Q�a�3>q��:T�:�HlÒĴ�s�F�ǿN�j_KB��j����Y�򕓅�F��m��y�������ә�mn2�&�^Vg���iA��v0'���5�:�}?J�u;;�d �+w����g����"��3�F�	}c�G@)����⩚�D�<xD������Kq>*���]�sq��ԯt@���������g�ҫ՜�3�ĸ<�����O:1S��&�=�ϔ��Q ��RX�#�A�04�u~n�!B��h�C	��KJ���?~�ꘐ&W�+eIIYc�g�Iꞕ#�c�~���6z���	^���P'�9�>��P��ڳ��.��u��K��QM@�Ǹ?�H{���.�n��X�L�=�orN�p�$��|�G4ˏPB�r,kZj�����.K�w"ߒT�����q0݌��q�#��-�yQ�:�e��'�0�Bu����|?����0��QK�҈Jx$�_�˞�O��p���t�as�+��J~���)3�c��)�m(�����K"eALM�Hx�+O ��5p���,�"L�1�󯏾�C�<dK�!f!O�IvK�3pa�����Ƙu#(�R�X^�ĵ�[[τ�o�֯�ܶ��vЉ���-���}�ȶ#~>u��r#P IeEzO�?���lk?]��"����X<�#�����h.p����j���o�.M��漱�r�7��6���^��>�;9�[|��J/n?�Qg�!隩�]�ֱEj��S�/�P�E��P�.S�e��Ǿ�(�$��%2���Y2�_i�����FXnr�m:��� ��x���W>��{	���g<WLud�M�X(���U�#窐SJ��ߚZa���A�5��|��A��2�[�"�[�b��r�����Ǽǵ�ٜ��DNU^��[�!Q}х��(�UF��~H�[�a���0�6��C��Û���EJʏ��E�u�͌]�8�h?�p*�~Ɇd�١Qa�d����bQ�٧(��A�.QI*�,tۣ�]Y#��bu��d�x�\����w�¤92F�z`��M!����0�r��J�*+_��>��y|����3��'���œ�Л&�}��:�]�0��3o�����x&1��q&u�(�������fUy�ϵ�r��m}c�Ͱ���ˡ�,n�@j�]�<����c��K�a+�o��� ����"'�����̥7Ҳwa�H��
w�o�x���М��lT��X�X�6�{Bnj��￤�h6f��*zwȑ���]K�9磽P���>h�֕w�����'4������L�L�g-� �7FÔ̓��~���d8`%&ۋ�%�-�ь��h�OL�H_�W���gLw_9����'��0�'H�U�|q�PO���U�sc%Ǎ�X����d"+9�\���9=���S��U�d�*�,��z5�xV���Ȳp���8W�=G:������=�R@���e5�d@���B@��R�!�
�O��kN��Z��a�T\��k�}���\�⏬߄ej]}��`ɡd� B�w�L} W[I�4+p:�c_����Epeց��;�-g,��W�<-r����y2b?{	o��Gi+}VNԄ��t����٬�J��@~�9>�ņ6hO[��sYIٜ������tu+,���18��a��q �O��0�O�;�e�Ͼs�8i�J�����Īm�ԙ;Gq\�S.��
h��PE��!��s��b��؅C��e���(�V���^z����e<�՜�<��^M,���߀�����G���i!8�;��>-�C��Cf\<�&����T�_�h0Z��)h��8�⾯��8�e9'U�`c������a<%�9�" Qf�����!n`���;�Ke�l"���d(�OS���qji(�[��]��A5�d&����}}HI)y��`�̋�*�6w��h!{c���4�Y'�2,��D�5���U��ɰ��`��U���"2,8I�dRu7n���j�ɽD>$ �w���90�H��=���͍� v�"��FdӫnU0��k�H�&~5���u?e�=���z:�Pie9��I����F��鿮䨻����R� �"-Q�4�����ˆ�>��O��Lc����b�$|%X�o��0�E݅�ֱ�t���	��*@aU{�%��/�?y3�ޭM�����z�N�e�����Ғ��C���[�p���ӎI���I�^i�_�*���B3���0��>��d��W�R��}�n0�0�U���Ġ$�V�	��@��Eq���2~������R4�����x����E�F�����0��wT9�/�eٿ4i��@V�C��Ӷ�J%ݑ�B�5a�gM�^%BW"6�um"��9rUfX r~���7)� Z���_���7�W�����}�4:�˾Ա��������U��wr���z?�Z4���SZ�si}qǢ��>t���d�i(����f��4��Q5%p{V٪2����A����X��8�ed(����U�/��jNO�d����iE�ߖ?d���K�rɎ�:S�`������<`������uK��G����h��-L��fP�ǔ6˸o��m�t!@XlxVHYEB    c397    2030���Ia���ف��Ϯ�A��~�g^]:T���6��\��ѱit�}_�wC2	YL��l.�p��_��*bif�� �+iJ�I.�=�	y@Of�Y[ԫei���>bY��+W��7�)�I����b~�֎��~a��F0e�o�\������������n�ң<l(�Q́R�����+��u*�I"����g�- >q�y�PTl(\:r^�r�t	�V=�,Y���@�yXټɊ�a+��|�����G�}�}~L��Y �}�pM=D�`f~���}�� ���W�1�w�����p�y=�$�x��G>`��`bu�;�~���漏�,~[qlUbj��}�����R-��C�Sa�Bv��D���f3�>�>��,
j_A�SY4|ym��|`|A}dz���b<0b�C���1��B��RS<�"	V1A���2=
f�������J�&zD�w�}���4t����2D�Q��Ө�""{��᫣(L���Pn��'��A�!����;���ŸB��
�z���Y��Ih����.3������J[�{K����ۭ/I��u�e?�[>��������c��B���qcu��}�;A��C��(C&k���P/�9�8>J��})�k����gCIQ�	��<�o9F�3L�2����]�\�R�LTm*�v��с	<����w�:s�08���6Z�蹶�xQ�R���Mhw�(U���ST�<�6��L�\�����C���A0�����L�g?T�c��
O��²���l�P��6�';H��`�ʪ$�
�J|��=o���������1�;{iO�v�3T�Z����	ˊg���nO���⇑�4sg�_"X^U�|�z�=���(�����Т�� 
����&����yv\.}�orL�A��hm�qk��d3P�1��ۄmMe���`"�'��d�y	�s��RЕ<��Q���R%��J�\<a�Z�ɫ.�So����2�6�& W���b�M���#�" JQF�Fl#N�`X<��?�c�Gn��FX*n�^y��>Ͻ����U��.ҋE��@�ʵ�K*��Uk���ʝ݈���h�6��Kg��� ��٦���*E�}G�^�a�׍�Ϋ��7��]wqs����:��w?CA��Ƹ��A�J�EX�|	�wW�=�=t��o�^�2Z7�"ӑ�ю��L��I�l��7zt�U����H�v0�~��뭭�2��2�������D�>�c?�?V�zgRͭ%�?�E!�=�{�$�ǧ��3�vQ��n�p�����2��&L��P���g�-o�k��px�k�����C��2TUO.d��2`55�]�t~ĞK�����,�-Hx1ґ���)ZMsմBmz�����d�w;Q���1�Q�X�<*ގ�T$g:�9����p��_�}�!t�~z��g�?������Q��>�M�����b��R2v�p��8����/tPт�����01&B�L�٪�dfȡ)ȶ*+�S�I<�;�O���.��}l��V�˕C&r���Ây	�r�Bͮ���Y}�Ccz��Q�OD�b3?u&|34}�5��X���b�"��:��6��_�R�����]�ْ�ml�]���jy;��8�_��f�ƌJ4��H^U�[V��Jqa��Ø(Z{�q�>�B�+��"t�y�Q�������-���
��=�<c1��;ͬ5��ڧJ>u�3Yf���\��GUY����n���w*x��W
@�X���]�R[�޶_�
q����[�#5�Qͻw�j�����bI�&��?S��]��鄴�Yz<�����Yl@	G�������B3�x������w��R�����3�x~K���?�'t���Dd�*�i� g�L�\�ի�����_�bc�8����7��Q2z�#>.�	�N���xz�Qi�d@K*ۭ]�C���;ԝ� )���"O!���~��ʹդ��[\+�.�v�>�KA�p:��&\��R̎��~~���9b�&.�[�`zQ/;�R�,P�9��h�b����0IX���S	WӉr�>�6�Ԋ	>������! ��^0��ev��Bl������Oz=,��z��ID��mr���۴�AX5ԧ/�>���FAo7#����c��}��NQ%`����� }��?��	{ch�	�I5���UG�Dd֡��Y2���w:-Vw���W�	�!i��Xi��JB$[)G�1mr�p����#b��Z�C͚䘊���R��L=���4��ЁWp�B�Ԏ�L�kQ�]>C�(ɜ ApqR|��!VN9��Ɵ}%��� �6�����r�!��������5�Pb�n��=V[R>�6��?Аy?��r�����6�5<C۱7> ��"��.�N�Y�d˟(G l�#l��u��O�C0��4ȹ�@Z8UeglU��ت��Mb��H�o"��H&4�ʪc&���O]� ¾���O_{�[C�xk����IØ��G�[4*_C����X��Q(�_ ��_+�'���lɓ�f��F�R���,s?E�r�Q��6�ml����ڸψ��H�����s��6�3J`43qm�H�ĝ'-��n��Pe�Z�S@�s�m�g��JM��&y�����֕J�C����m��p�m�����j_���B���5χ�\I������{l�NO|�mWz��a�ð��j9��_/�5i�{�+t�C��W�N�_���!�?��d+�r��T��˭&1�����eQ��y���L�
�Qˬ8�10d��j�fGy�(�Y{��ڑ�U)_� �f�ٌ�Do�P(X�uڀHoC����Y
� �|�os�m�NjzZ������ɕ��5W��h".=���v~)�V': � �Iɏd����pS����0�B[*-C�xdK�1K<�#�K��/�j: �h�(�a���-6��Yf}b�![^�3]�����ԯ�k�-���� �S%tU����e�78\��b���B��\�;h��:]��:�((���!�e�#}ګ7ܘ�5�O�.�6qDKbfK��f�7쩮.�5�	���fr�b��5b0J��e~���"� �NS�fKnbfA2-$�D��hq�<�!.s�n)3\Z(�p4�$< �����]�������5n쨼�>͓���=��6φ�8�z��W�گjp ��Ҕ��=Ă��v�(�JͰp{sKZ�Uĺ�٬y�[���"u(Y�Q���^���F���懒q�)�n>�`����x���HF}��1j!��Gr���Ge�?����oc�!{8ahR�
o��$9j;H8�b�bS2���F��h�x�/*�s4"$���N���o��Ƹ��h�=��5��T�]�ϩRI�������`Ͷ�}�l���t��7b ��,9�n}��.�?�ſ	�*�cG(p��˧0{l��h����Y�|��X���fs�U=��Χg�� ���
�˰���@h�	��n��hʌR����',-6�S�+>!%Ȅ��7��%?��Af/!����3�D��>�şɖv�9d�yP�!m��z���'6�I�NٺD�X���/$n�#��O!�g$"��BP��D����wC���3l�� �WCc���~���Fy���	uhܭϿQB$⫚`�+FÙd�\���I�uN|���Dh�T�2��
 ���ת��+��4���Y�T��X�蟱��n;>)����H���i�+O�'3��7�(͘=w�A��`k�l��_w/y��Q����"a���L�/��8W�)NGQ���8�[i2O S�X~�xf���� GR'*��=��������Mr�G�@ ��˨��&ڮ��F����Au\)y�U��"�f�
�$f��|�32�9� ���X�J�|�BiA��c���I������m�K����,��P���g�	%�>��I�P�~=8�EX��"F��y ZF�S�R�G!����59͙`����k����,�38����u-/���]�����[��Ǌ��/��,2E�3d��0s�rP��������`�7g�dCt}J+�gv��3]8�|�(��Ƀ�=��K;q���M���k���C�ڙ��R.�<�W����z�a^��R7�".�� ���3�����bxjQ�J�*���y}i�ƃ�ܽ�xrNj���N���l�~�����A��)=�3�2��o�̐��d\"P%���b�T�f��s.�*/�p�td���0VQC^�(@����"�ESI��k���6��xe'<3ˬ�I+?�3�3�T���8���|ڦ�!<��J��� �^DDЅ�R?�-+�J���~�,��p���"������o��C���u�X5�hU� ��\z8U��K���=����WU�Xg���4���j��Ӿ��_{V΃Ƅ���Z6��1���,�n���Wv��xz���l'��/��l� 2F�[	��P���m�jǱ#����GW�o��R<���~\���_���!�K�u��>���#��������Ҕ~ ���g:v���Y!��۞k��i���qw񍄯��[�0�ntX�>My��ߍ����_؁��|$�?�K �L��m��L����f��Qh���d秈f�E�1<�G��Y�M�lg3��sJ���F��ː\�s���^��G�&�6���w��yZǴ��vf%�ܲ���2ݕ�b������ Xe�j5�yX��f��Pmѯ�E�W��E��8���R	L^�3n�}�o�������S�p[!���I�y��:�</����7���c#ٴ�B6���0��?f�'ҟ�_O��c�.RC;%�_e
�~�����C�sB�.fO�,�������{��2�͢�d';a�����/��)����9s��Ʈ�f�����������X��N5�7yj�к�����U0Y�ㆬ��o��n�ְ&^]l �˭��Y��MC�%��-��dԤ|�5
�=�B �y��9I� �'>ɾ�[6� 5D�)խ�K�[g�F�C�Jq�L)Qu8�y&���^b�̖.�V��6`qn��"��E)�fʊ�AF�3a�<��A\(�r�^�[<�C����9ʄ	"1.և���s����+H�a<"��%
lt�h����eKѸ�Sw��Yh?)�����#k�����.��!��Jr��w����$:'�����fӿ�7K��^�A�JL��&'�	h�.1��� ��Y����E~���N(^��O�{�V\��{E�gu���	�mz?�uUAA�0O��)�ߪ�q�굒j[6W��/�A�>��Q�B��<�!��wt3a��9�)�M��Y-�$T�3IM��%�\�A?��~q�n���=�fΏq��� �)�0��~�,X��m��ظ#�䷛��ڈ�d�n���_=���ɟ��3��B�G����9{���[���I�AsK�xS_ ���+C�/j����n��z��#k���@]��kL��=(°���|!�����m֡­ؗ?�ZE��%�+B_� H�H$h\v�����#��o�,`�aı�)�	��C��[�նq;��3hPV���pa�jfJ̢w��_�]��$e���j�h��Lm�~��.Y�p�������^�(���\�״�.jy�Q�����6D�Y�+�'GSϔD��T_e�S-��m�uW�	ƯK"���_c�ܹ�I%�U��đZMް�)k�ues��%�y�3��+�*Bi{&���)?m#7�>\�r�5.��P`�^��z
tc���Pm'"l�NdĔ��oK�a�g����E�3$�\;��������s|�R�G�-(����9d�{�j�P��X�����t�>Eg�.1�]g�G=ܥ�G�:N�io�V�.�rW�Q��N)<𯙧!�?i�a�}�j��·�e��ٮN��Gl1�J��o�?j(ѩ�]��?����y��?�}�!ͪ���M���B�KT�؛{C%XƮ�g�RB�T�H>�ʬ�g-��$>h�ݨG�:^M�=���
�o{mf��"5(Cwb=����g�9I� �B�����3�N��X>'e�����7��T�R3C>z8e��I؇`����d^�({��f�VU�C*#�1�C�vV�U��ܢ��øk��X�+�9����ɯ<q�\�fk2|X�_""^"���I�5J�+������eI��j<���em�j�B�o[�ȥ�d��������H"#q0�_�$?*Iek^�cy�xր�V�0@R�q�VRf��G0�4�;Ͳ�+戻������ֵ2�V�i�紹
�Z����	�Lb��l�e�O�B5�V=3.�@EL��iF�{�/iD����CI�S<���$�ƌ���7�$���ZV���{1��z��b�dV`��[W�̿9�"����)0�@j��5�^vt��?p�I~��`-ص��Bu�C��~�J��I�Q<}^��x��	��/�jqFa��=�%̳�Y�Vg�e2õ>B
�V����RU�ᾀukvf%�7�l@�M[�U�1��C�V)�7�fo�N ���ۧ�q7�o�+�@���ؐ�_M����.��ɡM,u���� ,�_�a�ZN���S2E��6��.������-Rn8���#ʹ��җI�q���A��u�s�z3���5^PbA�琢�����c�XS~�h�qJJ����	]�l!�s�p� -8���7t���xɎ.f�>�d�%W�0�j`䕔�p���U�:���5w�Vm���f��1���f��4��tN����׉ySK��e��yC䦓t)Ջ��.�]��@-	A)�����lA+� �$+�|���hU�3�5`�)�yr]~T�XK��U�^�6ZWh�j���w��A&˂��J�]� ��[	����/2��"6V��?���<�<���ф�
�r�A�rR5������.�ә8J�:�V}1�O�l�Z?vq�ށ"gH����U@h���������;����N���W,� �kl�+����N�T�/�?+z>�]*�CѼP|�ۨ�'c��/�"�I(���Qs���9����ɓ�qO⛦�(e���zNZ~�n+�34�����Z�w�����v��E*�<���D��z�N��A�ȃB}6��z�s�ۆ���Y�,�bB.�n�FT\�@��E�K{���xB|┼���G=�X(�n�w��\����͋a>��\h?��ɘG��9n������[��[�2������m�0.07#}�EYb�\kl���,.r��9n�a���-#'���c{��V֜����|�V>��iOD��-j���B$t��؟���PX+S���X0|u�r�-��GgA!���,�4�T�=͛�&���s��B ���&-)Al��y|��V�s*R�#4�QI�5����ؑ�n!� &��S�s��fҜ��St�Q|�T�y2}wD�����"W�z�>�����\�DO�c��1�D�6[�޹U���1��֢n�ޯ�+�^ {z𑓱"����z>>���P�����&r�]�F#V��-i�]πM� ��K�u@�ZM�Jd�j�;�w���>��w2k���5Z�X�M�.(�H�[v��P~��jũr�{�a�d3�3Ķ����UV')W�Ё
;��/-�����Ǖ1��,|�o�n]���^��c�wͧ,-� �"� Z)Yia�+���oQf�m41�X�rc�A�Ӷ�N行�Lc��<W�80S����'�����в���&$V��O�~jD|,�( �mL�K��a�k �18W�d�T�y��WC�ߝo��"���ؙj���[H��ы��,8�È�y�6X��#C �4~*��C/��E����՚C�p�^�BL-9��*�s#�>�����7(�O��!Ǹ0OH��hH��ጝ282a�j.}n%6��{A��Am�H��"/鼶w�$[�-��6��T��Z�ܟ���/� �Ɣܔ�0��ҕZ���k@��_��y�l\������l�M�*�wjH��\��B*�e����dW�	o�H�˶q��RV��u,�'�=Z��^uW��ݥB4�/-����~�'��V��)���A��Irx	2!}�`3�#V��o�2�ܷ�Mq��y�(���
f#�/�r\L�����G���^O�c_M�zI���D