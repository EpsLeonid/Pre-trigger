XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���5��.F�K���d;��0u�m���E�]rfJ�����H۫`��F.Po=Xs�}��})b
T��n0��Z|�`I����[��3�2'���%e6����4�^�&2��c�.��6ȚX���щ c����(\wx���u ��3�CőL:	AW\WR]�$ ����$V3���������Pt��M2�%v�@����5�U%:cxЍ6��}4�j���-Ƥgq��c{�,ӰyF�-�!�R�3p�f£�58�.T�?]��B�n-�.��L)��U|V�q��պ�[sj0�A/�����f�cw361:)y�ZG�Qm��E�6�r�ςs��E7�V�"P#"c��anl��6�4$yq��� 9�E���n�*�9�Hp�ut�W���ܝ|y���~~�Ve'){ֽ�9�-�3X�+���ɠk`^��>���z6�����
��7�ŭ�ߤ���j62���`�ɬ�y�}i�H��:\��lE$P�bg$�pjs��H'�8�c[���[1���i��*�/���A`�GYi ��9g���dTK�SF̪���I�Ȱ�Ut�L���!ϲk^�xW)�����F��^���С��b�(	s˶O��9�T��?���!��}Q΋>�P�x�X��<�yO�� ��朼�Fp˟=��-���7��f,jJ-��N�2��K���}�_!5�H�-l*_`������F�h���yY~��r�^��()zc:dػ;��nС���P�<��^�'BT�-/[XlxVHYEB    fa00    2620n;�L�}��B��6S��sT�Ē������p�s��g�zI_H��.3L(_(٧�'�r��c!b�͗�UJ��,�ў��K�7b��:�.;���k��.�1=[~1�~�|��	�F����as����/�~���X8�ӣ#�Τ}�rEu��6^Ņ�#f������DB#v�N�r\�ݔ�8�Ň�a��G�R��W륡����\q<�_OolX�L.)J��ߋ5r�{(��	=�t�kX��2�Ɯ�Z�4�s�5&��A��3�~�m��h^�ٯ��*m*�Z��C����
�(^� ��6��ҳ3Ce,q]��_�W7���c5r��.ʐ�����	_��+��0h�H��!7�m��0�+�V��rN⯻|\�2���\,�ɰ�?A3P6�χr���Ä�OzJH�'xٸE��X�8>�t���-�o�%5�Lޙ^V9T�5n�G�|�On�@z�ozr L�����TN���O���Eb!|7�v�� ���ރ��#�Q:�}Q� �1���t��M�����-�-y,io�:߶3F+��Sv�2L�ʋ`D��L鬙�x0��>��z
���S����形�M%3]�͎	S�X�"�+�%ks�%FL7��5��gZ�w<#��]�D!Xu�*��A	n���+Z0�(�|��pX�4sd��P���MUn�e��<b��=ޔ�/�^�"!':4Ohc����l�O�u0����eX����qїq%�pq�a��f�h�}��.�*���~?s������Sx���+w��Ȥ|S�b��� ����;�XDVo�F�S��+8P=��0��?�W�^��4�n8�:#ϸ.0|�*����M(_*&��N��x�^/?�mf�Y�/.�d�5 S��Z��ր��9���al�)����#�F�C�VvD1��&&U&�J��K*ô�"),���zQ[�6N.�$�#0����!��n}n�ߒ�ұ�4X⃭�ܑ��i��nn2��"!����<��|͖R�b�;�Iގr"ǝ|cSnU�)�=w�dW8����l�Y�/�t]��z��DjJ۽�Ͱu _�0��d e[0Cq����a|�-a�R�S���ʗm�E��&�"���L1Q"�V�]���jR����
��_;Q�v(g#�����aV�)�v!t-�*���c��т'[��v��t�+�`́2#�fV�8@���*��Nh��FaqpǬ#�Z�<U;�0��u��|����\ {�T�ʡ�w��`?��s>���_�q��9�{��`�A�y����S��?�/r�Y�)=]I2 �m̓�		^�G��zg�C`��җ�� ��Ø�G�d\�^�SI��_`�x�n(���&v�s~ˍ6&���ި�����~�c'g�o����̩�G�ǀ/��}��5�`#p�T�W$"0�]��S�О�@��]�ƒlU�(N�>��y(;�1�6S@�݃~Z3������l��c��*���#"���j�-��a���a�_��z1��5��N��
��=)宮�-�ױ��p�ǐYY�ɇ������7��.Hg�2���gU.)}OY!���<���v�Ü�a����=K��x�o�6��9i.�5��j��B�s�ݪ�C�Hf�~��נ�X���&�f�9�|�*?�1xg)on��޳�-9O��4&����o"���DcSE^�/��Y9No禍c)���"�30�\�A-Q]�&�Rw9�e�EI�����K#�'�B*���%��Or��GV�WkQ?|�G�CN��� �0/Z�jj�D"H8���%C����%P��6�n�Ȗ��z��):����K���;���ż������C��lS!?@����GNl��e<p������z���ɃY+?�0�����{�Ib@6����~���q�:3Z�[!���jjX����Q���c����s�9�-E�b��]Q�? �-U	�oghgM�uM �D���F�QX���q-m�̣��ow-��7�*��25���غ?��hi�����������OkO��$*��N���<��D��f�n
,��"�v+���7Z���P9/��o�\�6 ��F��b��
j�
ڵ��'�.���!'�5b\��o�g�L������ԓ�̈����[l�J�-��F&�L�rĴ%�i��E�фM��Z���2�K(��vǯ��!Lɒž�'�Ӈ�(�aݯ��L�_�Krs�EX�-��0~��)��h�U]�I�F��fol92�?W��Ñ�͞����Tj�2x�P���55���Z�;5y~XT��Ӛ|�Ϩ��H��G���O6>I�T!U�����YA�/�`���;~�8u�E��W��	��)�Vv��Z�C
�ȀS�����e�:�)`�6'p��M��1%��U {�{�;'�uZZ|:Yg�=����ڤ=�����q�c(�z��e�u����e����;ƿ�Y7����z;|*i��[���ڔ�SV�Cش��}{���7W�C��k����h�vi������a�(��n��c���S��f�>��FHT2\"0,�G[K��^���Q�vӐv4���	QC���Z�dJO�<8��K�%ٚ��?[�d��<D36�Ad=����0i	�a�QR9��D��Q��4�}{Sfjy�jw�ˬ+9K��h�.�׉:��ߪq"��Zc���~2�M!���~�Ŕ�5��U}d����5v���r��"S���V�sZN�p�\�2R�iA0(`y�Yv9 Y��<����(ψQ9JB�'���0�'-�O�������mX"`�:�=�[g�	�rŜ���m�"A�8�O�i��*�?�n[`\]�"�5c����\�KѫPT�ԫM=5,��a����0�;����zl����ڢ�NT��:Ok~�A��7S�Ye�X�#Yb0��n��<��!;"r�aP�ۡ�]2�@�w;�<U&���ѷh����N�MA_�X�5iH���
�fBu�Cx�~��U�O&�9)��·��g�e���|T�wL�E��t��fbY���m>��t����W2�\�g�	��Ö���,�ar�G������#�Ԡ߬n9������D��/��9�`Ny8�|�#��5�cYnV4��c�+Sى�۵��є萟�~�S���Gz�ռ�W��kGp6�mf"�W�&+-�+|�$<ኵ��G{��\X��d�鲋�TU�Dw�5��b8��\|�]�t�H^u��7w�yqaK��?�W�^箞%�	$Vӵ%;D�� �:j�R��#2�:�d_i�]Or��5�[��Y���7@�~����z����WiU)�v7�����"�v�����1�1�5zD����.�%�;�p��Ƈr��0�a������٣!������>�ز��~_�,���)2����Ѭͼ�xzJO#�î��}�,g��[��5/8B~�,��MM��`���X0���,�=�.{�R�`4�_^���K�4Kj|B��ʙ����#�z��}��l$C�p��evJ�@QF�:Ç�o1�5�(�E��ϓ���Uz|��99�Y���,-Z���G�"x��Su뫩0&��-�pg^-�~��=ٽ=�T���W:�_��ӵ7�'���a��1-��*<� �4��;���K����gA������S�3�lC�R��"�N��Qi{��hw�jn7ЈҐ�Zq�����+��Oz%���?�Fo �� Q�4[�������.�?�ҟ�W /�� 2�^�_T��c�>�R��	��\Ƒ)�����K9�A�md �u|�>w{�o�('!��p `$Շ��w�����L��o�gܜ@�<L��o��:�"�0t���p�DeC�R[�*֣A�z��`�^�J>��h���Q��L� �@�{����滗]i�f$���eZH"�4V���Vh��ų�� �B���zL͛	U��a�-ٯ��Ugݺ��#d\%��$�@�n����A�B�H�8H�2m�ȓ#����,rv�Za����m����յ�t�|R;�v�OQ��X�hNF���M�5+��N�
�F���_��Ky��~w��IW����d�Q)~��`��ˀ���B{4y�VR�G�+��O��,�:5q��R�tj!�Щ���k�s_K,+9�o��������#^��vW�a����g�QÑKi/ �K���;t�������l�Z߄�Y��w�ҖOp�-"7���֙ٯ�:��빉�<,`�鐠���:�d����U��a�Jٹ�\|+�Qn7&1�?/!�e)�����n,Ʉ�O�u3/��
����9�<���O�z���ag�-1��w13������`�/��"���V{�u��W���*����:^��Q[\�D^���������t�������6�v������m��jz�p����:���Drf6t�s+f4�γ�i��]Y,����K��������l���k�+�7̲\�̓kmOI�	dJ"�U��"r	R?��0T9�����n����ui���/����x\��ذ�G堠{Ձ�,y���{��P @n)�̍�d�xx��*ϊ2��>�V� �-o�2AU���ޡ�u+�L��Ig|�VK�Rx��MR5Z��I㠢�w����+_�c����u�sw|o���Y�E����Լ�8����BY�Р�R_�� ^쥍g�q��I��X9��S�W1
T4��/���JHcd&��ӁU�%%*ku���&������h��pT%|u 1�^?u�^�쇑X�s�c���:���%G����m1�^'LS��iHC<�rV3�a�x�A�YG�󽷈��W�qb��ц:.���i-�U��? �FSx������{"���=Qm���PX��ˤ�8����}隮$,���F�Y���A7BL�E���T��^�K�v�V�nYKT�큾V�I��i�7�;k�5�6�x3Vt���*�Hc�Ӭ@c}�a��������{>��ql@�9"V�¿����pM{�I߅S[�ym9Д�%�{��!�p��FNϷ�JL5��tS�>�p��Z���wD���@ѓ�`b:���0N��D��/R��)#hx�4
�����t{=:c��b��hߝ�YF�(��2B
攸�|r�x�{P^v;�8)�ف�f���ڹ+2�4��d�v�ߔ�Һ1+r?v"���'�vm�̋��֝�����Ak� GY�e�;u
8�@����>�,�]T��xuMF���������͎I�E)`��I_9�ƶ�7�("ٵ��u�RA�Bʺ1�*��}S��)��Jg�68��"���LOUg���k�K>��Tv$��r���!/�A�(@ebΞ˔�԰ �d:�p���2�i=P��aѢ]|��/LiZkFZ���F�(.��	l�	+>�<3�0�� Ƅ������{��5���(μu��]0�X�4��f���9�����.W�?)�7Q(O�G�{�
��D�P1l2�|�a���3*���FJ;���s����L:l���h�[y�(?G��s��XP�	�L
�JI[���T`1��� �r�F��h�4�Xe ,���8�#q5�@�
�S�_�4�dr,oK��D�Dծ5��cC�h�[t�����Fx��f2�MA�t/0X��_�7Q�T�?o��V%�C5H~4���Eɣ�� 
z+�O(�_����T��?%Ih�<��T�ֱ�}���1��6m}��N",��=��)�"	�Շn��Y,�CE}��/��'1��M-h�փw�6ǫ�I>,q�s6~��>�иl��K��[מ/�����Aі5�^�a0%������-G�웷|"�5y�z!�^U@���bD��'`E3n�EuQeI�Һ"x tH&�|ֳ����a�h@�H `�+N��&��G��S�ֹ|���r��p���)e�%�a����]WԴ'=�})��Y��2y��wY��LG�$y�-�;�E�I���9��HiF��"�˳��Q
㣉U��As�B��T��Y�����i�o�6�gІ��i���ʅ��������*o�X���ftp�#�A��KJ9p�ۨ�,�d�v��wԎq�K7�H�����G�3ܫ��x��2Ƥ�P6����\D^��$�#t�k>>1V��G�6�m�FW���k� u%噈7����@��kW0/a��;��W���2��mv�4C�j��,�r�m�tɰ�)��/��0l�ȭ����'�'i\�Me��y�m:N e��i�z{O�/G��j�!��ѱP�|�j�Y��&	س��1n���gP�TQ?�z	f�m,D��G0�F4��	rՕl���&�Q"{�*�����X#䄮�C��"�'��"l���V��x�`"n�g}6w�c�o���Q0V��O6&Jr���~c�t�F����P�ZK�M��F�����5.�8z�KY�IUU�)��T| �e��l��Ou-����ś���ޔHˀ�۴���'�ek��e#�E�`	�76[��w������+�	@L�,kH���v�p�E@��NP��?P<�wIWyy#S����N�p���}R�9̘=M�fM��E�;ߡ����J6{i%'N�C��4	 :T�H}�������,6����"�iA�F֌�;ȵϝ�-�J�zx���s,Mܪ�,��J* a�p�(����=��V�Ա�S����
��A,�ERx�� �^|�إ�������R?���U�r8�[J�i{����$��TQ��@k��>^TNF�?�B X�"C�,"�Wy
���
�OT؊���pUYy��2&Ŝi�ye"���P?��T)��RK*�"��?}����4,L�*��->���
����-{y����O��;�>�=�[p`�`��n�y�[3�z&�d6f�o�][}+�)�DȱЉO�cڣ�����`з���Ϥ�g!NT!_R�F2t� �%ώ��*�yر� �X�a��*�h'�Y)D���簜!�"+��Rs_���o�=� �N�T62ډ��x~�.{�Q ��7w8m4�4�y���{��&���"�l��M�a��k���m��jrH��p�J͙k��@2�)*ȶ����r�y�[�k.���Uq��E���[�'��<�ā��_ K<��W^�,��a&����l����N:$�dF�>U9��#����6��_nd����O�d�4�E ������3�{5�&�ra�=w�(#<����(�G��iN��!ޗ%��fQ�{�Zd�h[NQ�vr���V��E�u����\G�=�`��a~�� &}B�}�=2|�c�H���sA��U��L���?��������	2h���ؖ�ݜ_X��r���"�����1[E]I��&P��5��M��:�j��M���ܛ�*�]S	�DШ w�$w�|*]n�6����N���2t�j��8t��|���g?�����d�2�HY*�i�>J.�PU���+��{;7��e���T��`"��ߗ|"ўrT�b8,�G]f#!�����$3 j�=`���a�� ��������%朇���0ʞ]M�{�j��e�d�z<�����}{٘�M��Tp{�a{x����������`��������v�N��N2嬟�{��T�x��m�o�i��k�E*bs4Tb�zӣ����}�����iqL��T���?��"u"��ғ�nb x6ؼ+�Sמ"��v���9���N���g��X����/��S��	zp<��3OEI9�E[��>�zn�X��9ׯR������~�WY�m��K���Ȗ���ف�!������4�t8��P�'��*q�ː���S��HX�Ϳv����C%oٙ���@��Xg|��ϟ��?F�c��(���4ц�Q���)-!ߞRލ��q�1\kG�A�8}��Rx���ރ0���H�y}b��n|�xD��?����ļ!�Hڹ���Y�0^~�,���P�˧n��2�,9��O�J1)u�r��I��փzz�aT�W ��|V�Hi�R���v�Tg'8{`Y�	�f��ˋ��`��#T��0�K8A�/7�~�g��� �t@��+%&B�宣�4v����"e%#Kyo��mu��by�]f'i���8FH���(�̎t��فI���u���CO%���j��D� ƀyR��c�魞,���C������"�Ӿ�7`����uԺ�9�L\�'�i�⑆�=n�@�+d���(�/�E׭Au$P���q�����kW�4=1_��Z����9|��I�����m3��g�:�T�8&~qH�� ��Pc�����W�a#sxB
[B�&Weէw���(�+·*�+/h%w��X0J�ɞ��Ԛ�'��#�C4�e�J+s|���Ȋ3�d�K���k��X���-�{HM�,Q�f��J7������B&m��2W�f���?}�V�C�����tVĖ�� 0�ǉ�^_f���}�u���9 L��b
d����T-3����� 4����_���G��P�p����vH�{�n��S��&B
;�$�7Q�#-�ͨ�xe�,����S���3.�z�P�'5p)�h�������@��hj&���#�N6�-��'U����wo~�	W���!
i'�°�N�54����@�cg�@�w�0�r�{�)4a������udg���^r��ku��T�d%�HN��Q���1�"���]roW�<xXϭ��&xI��P�p���0�^T�F�8�ʬ�(G�f�� 1�~c�b[_*˳?7-�D(��ޔ�/ ���R'����s�2� �'S�|����A���������qCn<�H�����C4�G��/*ri���,?���B�C����CwI�k%H]u�����{��]r��>K<�3J��E���Q��3���P��g��͉^y�<��ϗ�?oV��zA��X81�X�4�$D��H��ځO߆�Б)�tx�^�d/����m�<�t������=���{U�}a�Ϟ+�P:ނ�����xZ�2s�r��G�EͳNIƘ�ܹo)F��,v�C���z��=\7#����-�M2a[��;q$�DٛY�p��F]�/�OXԹÐ�����J���g�"�JƠ�I"�=̵(�e��	0�4���0������;�₮�&\#d^b%�
��K�毘�1������n־�|b���:����V
��ki�Ј2d�b�Q��kv��� �.��H��ܘ�gL�/�Bx\{�����H��cf/��
�[�LV��&���Qw5��d��7�1�s�V ߵD�u*�����������.]^��i���r��VC����齆2/�I�P�w#�-���6(��w�>�s����Ƞ��:�Ψie��v�0L`��|�m��)�+�C�j��[�)��z����� �ƁB
#XT�g���B�J��<"&w���%O������EwW�0W$��B���\mK�����6�Ϧ;��r�r�/��&'G�^��m$����hxͶ�/i6���[�&��hu�/��=r�����MyR�|o1ƳU��5LT���Y*
;9['�M }��my���bi���h$����TJ�ǐXlxVHYEB    37e1     ba0�<+�z�^;K���KkD]v8�ufyt��0� �0c��mSe;�]��Sg�3ām��J�,�ztMpbEz��1�]\��a�$�aM"�rȩQ��=�v�6�mm���-��д�]8�`fY� J�GB���;�/ƅU��o&��(���_F�Z�U�P�a5��<��\�.b��Ka�\�[�n)�� ���]�{�2�/�����$�q������ˇ�kuP�H�_��\�k���qwL���E������K��R���V��%,*�L��"g��vLKK[�2�i`���Mel�q������JU�*���[����U�}��ӟa�d���:3/�8�b����(�v��p\t��~ħ��~z�ߓ�u�-i��9j;�K�	���~ *�)-��]�� ���9�O�g�C~y�feݘ�N������x9�ldDb7��[�d�%�?-P��jk~�0zB��Gq���0��Ņ��(��2M"[��A8��5߼p�ode-M��O�0���r���7W���
�(F`����2���;~�}�|:*�򖉱���%�]e����64��+6�*N�ȓ�cO�R�_�����;���ڕ	�6RA��'�����-��Psc�¸E����=ԧ��$�0�Sg��$)dq��A���-�r������X2?/p��x�y��R�;B��)ƙ#Z��=�������)pȾ%=�Z�z.�6�r�=n1hq;w�)/��d0jz��*(WP	|*)[Ն�K)�-���GX�'������Mx�,�\ z����ְ��rly��l"?�^�y+�,I�,�`3�}{-H�@�&�K��9(r��gp�xz��,�oP چ�l����{h�92��2�`��y##��yZ�p)N�l�st������%�����g��|���h�0��J#ACz����4-���Ȭb_>�o���oE���stw7o�*�,{�DqKD���n�����K���0Q�9sZ��MB�dn�{G{G��`�&R5U��D��z �S�,��_垻@Yљ���Z#�c��y�nr�)S������Q=�ڤ/r���8��;���di�T�"���|í\�����;>�PK�:� �i*���MBH�/qZ #%��Z�k_��շ��iE�������!(��7��#=2�9�b�|~�딜^dK9׿�k�
�,�c��H�����������w��`%�F��^�����&0�'�/��1޻=D:e��>��p����=Ǚ^Ԟ��8�:8�"��$R`���4�OJ}���\��C/y.O3nΪr�?�C�燮�E`	#��1���cxEjA�!�D�Ch�'*6x�̣���Kv���^�y%�w���W^$�8f�hzǪ�H�H-^rx�b�oG�Z�579�Rn�E�%�{��p�j���)z�����w�dz�c�::hn`n��G��թ�Ļ�im����^�-~x>�w���Xn�lvV�b@��4ѡo��-��Hן�ޠ��|�<�]ظ��L�!��_�\�ӧ�Eؾ���3�+�#|��_x�cԷ�r���E�b�_�(w_dW����'o����m Y��&p�	�2�o*x�P�9���{�{�G7�{�Ew�Pߛ��JftW��6�t��y�������v�l�7�?>1��͝_�N�K8��Qr�n)�9^�Ѿ'dB�G�8�,��k��V��?7�˭�Ak��.��H_�?�m�th��bB�� MK��!���V�f+G��,w��H�x*+sȝ�irc3Ŀ�����&]/�9����h�˷�4�qVh������k?A��6F������?��EvI�L���Y[p�-F���kv!jkur3o-�)k��|=�Ub���7{�������n[�e�dۄT���ؤ��=�r=ʎ*'� cʱ�"[%���{�Y�p�@�VԳ�2�7���qh��nV�SJ��=^k��tr���c��v|��J�	'R����P�l�Ʉ/3 r#u��zJ!+�4����3�m|g	�tCw�Z<*�;f!���P��x�8�w�PP�rK9�[V}��f�}�Dg��Y���P�ȪxnyHؠI{ l�T���0m�1������Q���~Y5{Q�x>�ڶ�0�1&��z�n�v��􈻯���1�e���I��</#!�k,D�
	e��+1�N'�x}����}�q@U$� 2��#�����2�$aa�PA��O���p�u{����^Y����e� � y@���Á��9�33���U�����j�ƕY-���32N&�l�LX�֘碻ma�mC*�U��d%�f�z?{T�]R��>a�B�hyp������
�='�$�Ea�1�[�t��*���XB�
�����`�6�}���Q���=��Mi,��6�s����+�"�z)����J:^A����	��4Y�ln��v���o}f;rf嬹�v0Ɗw<�(~�r9�YP�;ΟG�~r�Lo�Z�6��㔇-��x�8ϐ�}1}��e+f})���x8A7��>��'Ue�"I��TdW#�D(Ʉ^ו�b�ݶW|S��=����I���P<Fa"���޴��0�oW��(l`j��#�}/��"XY�$<��U�h��`�7���EY3��i����Y�{!�%8O� �<T�b�M�m��v�e�1y}ؖ �
$q{dB��S�K��v+��8�'��0�=4�?��瓲�;��%2��%$eREP�n$�Q�6ۆ�r�:�M?���l���-��L����)����;n!r"�i���5c���h�3Vf2v31�[ܩ��.Bj��8��'پ��j����s\���9�C]|��n6,��T��"*C��CT��7�zl�@N`u�v*�*�cd��$�t���/}���� Fp{�k��r�?g�f��