XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����M��SIKY��ڗF���$�a�nv�(]˃'�a��0��1�M��Y/m��#�6ek�៉�@*B���9צ9��W��Iк\�%]�DÊ�^2��.U���,{��97�TVa���\2ؙs�7����OAYaq�*�A{;��g�II��!�u�*}`���3$�-�G���ipV��p����#��I�,E��`�Ҡ:XO��d�7���T"q�ԃ:��Q.��~�tٍ���/$06/�f��vqG����8�h�3��V�_�v;n5��¦��O��^��)0�lH/��BX?k(���=���jF~{5����c6������dS"�i+K�\�5�=2�䂘�N�N\]��7��#i=dJ����Ѹ�� �RK�΀"3M8�^#�F�	���3a�����w5+���M�� d��Z@)I�M�IQ�:"Y�T����͜B������1����H|�*�LԶ�2-m��^KȔ́uὧ�D��y�/�s!��[υ�a�N��':��yH�(�_�-8hն2�\RԮ_���@���Bʳ�Eŕ�>�tC	�������8\�M �A�-�����wl$i} f� R
s���̦Z�'��r���0q�'#��'�YHM?�DLq<����-	�D�}Hd��ԃc��Ej��3���[�3��7͞'�$�i$�9W��#���_�9�@��u�!!u�M�k#ڔ�T�$����,�cR�[І�W>����F@Wt�6�VQwh�oPO��XlxVHYEB    4548    10a0R�+
^ÛVP��I-����S�Oqe=P*r�k�3�^[�:)�{z�q�}>��w�跄�=K�Yh�hjV�a>�u��D6::���]0T	"����(���D����m�r�����ki��)�?Nf˰eXO�^�2<tiܸi8��9�ݺ6k�`&�{� E��z��M��(���.`8�ۘ����M����uA���k'�1
dv��:J�/\�W'[�~����^ʎ~����)�PQ���<�`���i�w�����^!�џ��[�ľ�./���&�P��]�5�?��'�z�9+���;�3䪻���C 1�i�4]�V{�7�{i3�[��b�8Sͽ׽�[��N��Pr;7&�z^76ET3����׽��Ta	��e^�þ���|� &� �	}��CG'���8��큼�*�� ��}��r|�-�J"*:K�j��e�8�����Kx���ඏ��2���1ZY�Q�w�ܗ�.`�L��ٚ�w����r��]W��pE�RhL"	�@JO�I
 ��=�c�s�������c�r����S\K2 ���� �g"&��M�#� F�ļ;p�nG��`�m5�F�����C,�R�I˪����$����B�>V�шD�?�����t�S���	@I {��
�7��#�7:;ӓ+�_K�	���mߋ׆��WQ/�.��%�.q��c5h�HROf�����P?Ѷ �}�O������^����bp�.]VƗ9����X�J��+����Љ1 ���h���T������USq��XX~*�\7H�l�� ����j�i-i��*��M����J��ɚ�0�����yyމ-P��u5Y�޲�q^x�B�<6�J�F�mT��X?��`���<c�g�|�U�x%��R��	�%!��Ʒ�n?Ј�lk'6"DBGC��� ���0,�N>��GJ.�����:oJ��ΰ+e�?E=&Ս/�.߬[�x�ʮ̻���􋄻�S��%>��K`�ۤ�7��Cz�".���9�U#w^�=��r�i�����_�������BK��["����{��-!�e
�Y��px�#Zc=�����4��'�a�T�Bzz�0iVU�%- �]��!Q�~JC�)����)���	�L4�p���_HD~��d���I崽u����|�5�g��D�|~��Vno�F[K�[oh�S����r�!"	5��mAV��1�o�z�"��>��>p!,��y:_!��A{ofgl%���E�b�48Z1x�%�.搩[�� u�����a��c5~e�V�|R,��� �o[K�O=�Q���Ifw�5e����j�S�.4�b%.dcbM�{�&�oJĘ�����Ѕsz� �{�g���?��h^���wN_����[�Y"[�q�'g�g��#E�i<*e��9[izW�7�&�nH>_߮��������VM&���_���2���t�;����<���(������Z�i���L��:x�_xt�S�jO �$������e�<�Z�F��F�:�̲��:UV��ָ�� /B���='Y��Q�0�Cg���t
i\�-w�ãC����0[����8�#��<�l�uxǸm����ޘ��%�j�{�w���щyO����wJ2�6ɕ���,�����'cV��b�q�Z׶ْO��b_���:.�G�A�u]�Y'�z�x�	&�y��mK>��v��cT�4b�<�n2,�4�����P��d�h�2{�_�F�Hޡ��,��^�o؍�9м��b�4�u�,-��d�o��U�>K�Rj����P8?�g���VDc(Cz!:���Q��ksAIw��Lt�#7vM�e�G[�I*_pS���&bc.F����ƀO�� X-)�C����Å���BHl�JtP�Hߝ�Tݓ��i@�{��h��%Xy���0Yv�ql Q�����aR�LqRj�>ƍ�9��^�	���͡�c��V��XQ��T\�Iq�}I1��R��fu�f%�ًӈ^��Cւ>M������u���h��#�	�u�]9�n�68���z���:Z�\��龅{&���݄��/�L�A�4}��u ���?!X�/+,0?�r������Ҵ�X��,��8��d�cPQ���j�<�dӹ0*xS5�n�}�S��撨��['�l���lY%INP
cn^��>�f��=i�~,���Yxhk����L����'�8��O���ϧP'M9[���&��^t?`1��\��MP.1�[!֝�(�u�jb��Q����D�H��c.?ޤ���sH-(g�tV�`<>^���5�~��8[n��j|yX���f���(�(���+&�W;���\�<�;�B0[��ˠ����K&�Ʈ����E!�$J/�ЇK�3��SӍ�虲G�?�h����,�\��+K؋;�ᦖ��,����L]��*^��;��A�ߒ{)���dCNI���|\�|�L�ꂬ j�dV�|X�b��ZZ�yߤ��t�9�]S�u����As&Bq��2�9':�O��⡡h�פ�0�֔j�5H�� ����϶�'��,��Z&o\���vyH���^y�r*�a���ֆ��3-s�����Ŧ9N@6yWGՕ�	�7T}���uW��2J�{t�M�>�&Rhe���*�Y�kE�w���s(C;G�i�?�9��тZ�W��ؼ�U���5rJ�eSa8 cU��k=�%��E�G��
ʳ��W�D�=�V��`��{DH���\�7�{����&C��ix?��L{mU+�?ď�(�lFpXGP�ɻ�]cky���f_<�u�DU��a�g F4�X5'9�L9-�j!JB���2��plzz=AQv�[�
�"~`v�j�bVs���(�'S��`_�h9*����O~�O��K��� p�~А<tNcS<�t�~�a��1�����P�
�D�E0� :K�O�,ʿ@�0��1gL8JYj�菗�p>M�Go޹/�ح�B��{�a���sp������Y�iƵ8�;�8{OsA|λ/T���=ƴN<֓���0P!@��_
�R������x�+�?�O�#5O����^�X�d9�I���$ B����w�ir m#�?�~�I䞴̊y�,��洷W�L�T"�5�*G���-6?�lCV��D8�цfx	%����Ά7T@̀�k���{p�E�������$(BwQH$�g/ f����d�!8⃣5������r���!��_T��sh&j������t^qZu�O��=z-�1
ʨ��r%��\�Z�U)����F��i�!@���{n��K!@�W�6�"z��kU�'�s����!�OCD�O;ig��dݔZ8�6r����n>dC�R��"��,H�3י�������Hb�Eb�4䀕��Q}L�J(� �`�13t�D�#V�m�g�����׳w!A@���{5�F�-�a�]�L�Id��wq����,Y�M��ŌO���ַUQ�4�`]��V��#�YtS&�r��Fa����ԯ_�[��M�ɐ���bX�����vUw�#���-�����oNN�s{�EYA�p����*�,a�y wlh'Z/k�����DL;X����fJ�H�o�GZ��F��Mh��rС��zW�\�+��'@q;mY��p}��
�"����!V�D�d&-�x�o��g���V�H_!�n��l���s�5P^����8α���J��js�?�sH�Y��M�/�z(*ELq^Z����j��t�>�Ί5��v��M�,��ҬH�e��c�nZ�I��jz?jɱ+-��\�#%4*���}�� �I賩�l䈯�E��DWZ Bb�P%�p/�������A�&�܅���e�4�^$?�u��u��#"��*}��VPsj.��Z�����`+�,�H8�"�����1��E/�MW��TVԥ���ӳ��(ZV�6�'9���C4;=c!\C���[>��pZ��苿s_O-9+�o����0Ç+{9ݫ���C5C�B��i�S�T�7
���\kG��&�q($�n�����qDO]�}쭧4���3��-��>?1kbD�I�Uÿ'/{P�^ :y�s!��o4�)�6�

�<�1JH3����]���^���d��X��������|�� 6%Ov���Ƅ���x�f��]t�k������u3�81��y;��J��������