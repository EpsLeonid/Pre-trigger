XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����߆h��ԁ��P��f����GP4c�bk��$W�_��C@��+�/#^zN�#%3�E7ݮP��_;\4t�� m|81�.kZ���$�6��<�Zk��j.�7u~%��i�<3:�gܕm���[^Ak�&o�oE�!n�8�#*��hߎTws���� �ku.�B���y���6FG��&�Q��x�3�;�fެvX��=�XE7���W��W!
�� QV)݄t�9����0����;J���ڝ��S=�補��3ɕ7�Z&�P��-�Z#�q0�Yd�dj+���a�Ag�����q+x<�� [)�ߺڮ���q�E��
��;�������L�ˊb�m��DI�m-�|���-�`( ZI��`�"[�w"{x���Jγv�xV�~��o�|��B+jB�"�'��S0��Sњ����k�G�rMj��a΍m�<<&��
�#�76�U
{�w#BФ\������M�$�˃��<\G贈���R��'rt���F!Ԧ�( ��^9G���@�ZC8�^C�8�'^Bl�/�-��5o҈�f[�~s��k�ڀϦ����E.:#'`��R8	�5,�g�r��%%�޷�<f$�<���^�.���R�Nl��v������Rl����n��%h��?���G�����S��dx�: ��$��*1X��z�Mh	�͍Q]"�%<ٻL���gȓ%G!Pi��c�,����w�:{��6[�O���j)�8���rNB���z�&騙e�XlxVHYEB    4c95    1190���8��0��{�D=}<Y���[��ѷZ�>�7�(e�,���(����U4���C v tr1��虛�ˉ�y+M�\�^D'&$)�d���-��II�~h�ֆ v��,�PRɱ?�ǽ�f��Ĭ00;��OaX4_��S$�#8�ΚBi�o�Ah��Q���F\���zK�g� x\���y�*WV���!L��d:�a�B�۴2W��H��j��{��~>���+��l�4�V�S��/�5���/�����I_Oe���Q������lMa0S�ʖ��S{(n�7Tz	�%�DI�\D0�P�E�B'f�5���{��=I�)��y�6�#C~�g|;���z�L��7���ew�\BO&0{<:���6���M�����O�,�~ι@eX7�]h��X#q�"҉C��6|�ֆ��jY�6ҫ"dAᄄ�G���s�KnU�^8�9�n}�>���Ծ|:!m�\�7Y�'�R�d5:�P+���-�0�|.�a�BR�����R�H��﫱��̬4��O���T	�\�����og�E;�ͣ�i,��"�.�+q���e�����2�H% ���t��r�#q��v� ������&c	E��sXR7�O�U��5�F�I���V��q�+9��=�I��_�V</[֮�"=k�)w�'����\F0�AlKc\�%L��Ny������̴�4M�$- 3���� �(�D���X�X��u� mQv�^%�H�㟧R5P [���o��+B�u]�%_FR��bd��AZFɢg��)�'���V:�1����<3����i��k�1D���(����`#�-��;8 \T�G�U�|����n> �/P����9�ll:a�Y5��"�_ ���h��,�gi#�থ5F/�g�Y=�eYlz�@��0��d� �A����o#`�k%u�qx�ظttەd|m�U٨8zwW����˔��Y*4S�[G�I|`�f��]7�lW���u�6�:�Z�p�7���[�6;Hv� -��EQ:�=t�j���ҽźRTz2ܲ��8���C~�w��L�!���M��jٲ���O<����Q���*^���-{�(C�A�� ��J�Ti���$kY���Հ"d�+�GNl*|���T��Q�Pl�
������� ʃZ�o��%>��8O24���V����\F"��z%�mH�g��S�H�m�F��;���v��0d��H��D����>%�]��O<1Q����I,ٺ#�B��1 FQ_���x�N��L�����q;�1��{��߂��P�Q��X���k��w$YheUO�1���E��[��$�{�����
��5��\��v�3��=���ȱ�����P�����4�Z_@Qh�[�T��@�bްc$�"K�P
��Ϧ��\��,�T� �r��]� �4@XiZG�T��D���5J�Rs����|��> �l��&04�-7��"�q�X�?�1���H� �ʍ���H~�Š�Ά�*�C�ry@��51���V�fc��K"��B6TH�������S��}d0MVk���*\�{<�d06��맟Q7˻+�)_\M�oy~��;!#FnF���|�6S���5pn� J��X�Հ�1�|��G�MD)�k:�;�ۋ�5���(��?�,pb��*���_��F�t��Bp�
h���H �����Ƞ��D�7zoX#�IU�m����"~�Pُ}�Έ�yB ��²rz{e$r�MK��"[@Q�O8��5�6�#��9[�SS��p�!iC�eTWc7i�?g�7t�����d�#eic {}�m��t��W���.ad�&˾���mJgo@��6b��sJ�K|b�Fz(�Rx�4��ܫ�겭����>FF�ՠ`0��:��s���h\%���V��`|2*�7���*H����fu�"�힘&v:��h�*+��`��[��~R_�l���p�g-�~v���0�6�
���������������a�K�>�4!x�0�mBޘ����6˸�T_�9z� �!�q���~��	5P��C�?24I�e왜���[�y˧d����k��"MM��lP�����hLC�F��ѫ��8��9K_�ht�|uf=��b���qzP�>2=�5Kg�\���poW9л�����O'�T��ȨB��|R�¥(/��T�;��`�`ht5	�T��# TȬ,^=�����M����܎��[�J��=]Ρ��MQ�`&���g9�+�:�[�.����b����9R��oq!mc��%�nv񙶈���t�g��j~��:���25Q�qh�c�%�9���BA.�HAư�N�ط��q�DȢwȈ�z��j@� �i,!7�9�#��B_�&#R,[[��X\.�F��^{�7��!�Y����[f�I=�c�Iz��Y�����o�ºrU��DX��J�t���kS���=�[��B9n���&y������޽�헖�d[���:�+<i�A�x}Y�h�۹�1�pW�-���á�b��"����-ܩǥ+	��0]S=�"s��rc�K�
��B�����#r֢j��ܼu��������遧PQ�g ��(o�`���(��#��)a0��̹��%�T�!�5��p	�K��#y����UF]�N���`��c3U˝Lw��X�B�͵����@(P
�|�#jq�~Ώ��P��>Od9���D
{�&��+^o�g<}4D�*/��'� C9X�v8��;�ٞ��e[�u���y5�FW֤0*7y#�����m2�F��a9��� �@����<vm�1_d1苸f8A����/d|d4g�����⮬���U[����JJ^+���z�g�k)bb�$I�M��Z��p���5DC����lmp��!�F1L�cg�Ex��5���`���3L��v����MצŜR�3MһI��<a�@=Q��N�7�&��w�NNa����G��2�a�����U(W��ѳ!��,����I?�~�J�sPmvr&�r��Dl�w�ʼW��*�.�T����b�*� ���g�_%� �<8�9N�5�U�A�E��̛7�L�,G�2���V'C��˲���A���X_!Qa�K��l�^�h*����/�Ax�nAP�0� �k;-@�I��őBݯ� X�'݄׍/�Վ}V�8��`�[�T���~�R�y���Xyu �@O`�'�%x>�b�>��Q��=�׏*�`Ђ$b�H��T��h^4�:��]�c���z@,-�G������_��N�4��ZF��oULQ_(
�q?m�vk~�fD��"�h�R�ӕ�
�-n`��n�~|����T�C�����*����= ��&i��R���bg<ܥp��NrByH���
��π(�ٌ<��!gZ�e<4���a���I�<C��ׁ}Ş�P�qHu��(��x\�ȹ*�UFP>,QRQ�O[��LW���P�n��a6$��hH-���.�4[	��$G�,�Tڥb�����\�*��1��:�j�L
���0��Y�Of��{�]�A�}��D}��{��7;C��;H�]/w.�hj����B�rG8�k��%�u�,w4��ݺhe�"K���l��k|���������-l|�T�i���o��������1A�֭t�����߮tGc|L̋ϸ���?�K>u�X}=���ȝ�PI�VG$0���c��&0˥]�!4PF+��m������A!�I�-�5Rp��"ҏ�������� �]�K^�'A��irT���ߗ*g��!�f�C��W&�j���~X΂UT�]j��'�����/���(x�FjJh5�bU���2,j{��ؖai*S*N��GcN�-1fY���F�� �������c�S'y,��x�o�#�X=)^ۏ[�;cVѢXcVB�Gw)���D<W���(�gρ��L���O�y��h�cN%���@5F=�>;n��Ƭ% ���=��r�r��~7&rs���qz67�r��P�n4��'�g��uDėI�Yq���)�WGWu��@�ŗ�s�� 5�H��JU:s��b|HkZ�v�'.h%;-����Z��?%���F ��.�|�_a��&9�G�:�	C�%�b�Gi8�۾�6��|��<�6;T��J����bj^�uuT���Нb� �tX�(�ȩv��Q-k�� >�e����J�	� �Y ���C��@���91�e�E��%yk�A9�N���I���*����;��r3��O�U
���;��ь�1��@��	ڱN;R���S��qjg�y8���dD��u�^���?������\������=���z($Ȓ�aE���S��DX�I7�C
*�a�U����xAZ�!�5�s�'�㋩ژZ�(]ʽz�7�I�6��&�{��Q�;��[}�z