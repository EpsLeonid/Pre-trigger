XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���i��i�.�ͬԘfOp�*߈'�����c��u;�����g�N�k/��l���#뱛*Tl�[��p5�zF??4i�����-l���E�W�2�`����0ÕU#�qڧ4����!��c�����{&���@���,��F�b���/=��C��s�~�z=|� ��޳����Dę���e��m�s&9ýv�������.TP^���Ca�O/����L0�*�R�*_�p$7m����&`��s�b(��l}K�p�� �G]��ٷ�=�G��5ǢG�-CNc��عC�#�_�EM��E��u}x�5a��� � PĬ�@�`��W4~ɌoQ�k�v�P�;��+������$�d�6�YZ"�G�?��[?{�,#��.� ��_�9҅�?D7~�J����]����R������X92� <��A�Hk�8�P'�k.��up�؏J��%��j
�n�a�B|�k���������	�k|͖{z�2�ˌNn��k�%���ꉐ�P�����AE���0Ʒ'b��
�	X	�L���+�3\MW���E7+��x�1�$i��bP-
~O���OĚ_����QTÜ�����U��@׿�!4�_�M�Gi/I���'d�M���2���%�u�9e�������{�1�%�j�k����	�GP=t���auX�"��/ ���I��U�k2���$c��f��s?{7��]�`��z���
}�CZ���P��XlxVHYEB    1eda     880:.��� ���+�3��"��x^4��"��lr��7�&�݌��+Ʃ
)���k�ԕ׾�����潷����4 �����gY\Sv��m�'�C�«,�-�;���_�v׎[�XR�[b��x�-���� (�X�:���-��?ep�ɦ�3�xF����hW�=�� _��7�8l���?��ǴiQ���f�'26��_�m/]=<@	�Y ���هn�9����o�"mWv�Y�4�	�Ͱd�k�S��8꟨��eB��d|�r
��	����csa���4�BM��z���3W��%{��cU��Cy�	�ޘ��#h�>L�ô���T���ۛ|��:�����̓�1��*σ�Y�=�+�N�}y,���F;X4v#��xof�|[�d��,���E�y:�
�+�]@L����z#h�Q(z��PۜX�{�� ��g@��N"N����v��i� e��ɛ�@y����_v���] Ĩo�88�DJ��H�a>y�Q�����8ݹƮ� j�i�ln��;pr��i7l����Ǫ�uߗ@�`M���mq�YJ����G��jC�
��u�h�#�]}�{b�m�u�è��&��d���D��݆������s!ާ�̾������~ZL�����^Q�||	��|�s�}��J�&��kyu�Aw��g���-[/��F�e��hq���a�H�8�t�8��ZR��Fa^E�)�*�i��ke �\��*@1��Q �T�]��0�g-��>�tr�>� ���M�R�臌B"������Vj!v��K����Qv��)��K��w>��x��󲑿ƞUXI��n��%�Z �T[�H P��u�x�fh�;�i�k{Gw�'����Gꇱ/�y(�Cj8ֹؖQ��q�X�.
�.�҃됐���ԥ�7��LJn#u^W8��+�5[��&P�.���Zf�'T.};�w��ɭ�e��C��ɞ�8��o�	��%pK�����J���r��]��ƗK-j��Y�	���U\�Q�[��C,۹��!B��Ym��|���>1P�.uЯ:I���򁼰�J
�0L�c��dF��&���R������<�#R3Ī����1��W���Ȍ�#�w�ᗝՎc �߇�:��C.m���~{�^ZJ�7��� ۳Z�d�/̝SAX_��'�1��{��H��:�̮A�*��0���+Kbw<��3Ƞ|�}�4dy�2�_
����� +���E�V"�%`��H��ō8�������H���*��d>�\!��;��4K`	m��y�o��^�]�����f쌔�cQ"	��t<O�I���گ.���wEq���q�]�u_�:�>�a%�������FKwgP9f���n�4=���~s�}��3�l�h�z�� �|f��1��*<���s+��^�[͖��4z2"X��l�s��bA*#���i�6g���%����0�H�p��ru�(�ရ���)�p�<���4#5.��70�+�6N��AE]�*I;�����2�lK�&"i�I��^�c�±�I��@�H��Y�-.�v�h��m;���&�WPY�zPܡ��>���Q-��v�(Q[̛%I7u�N��8�mix��F���Yq��d���x�I������@<��^�O�ɨ�7o^���8�b*�R���
G�OY_.�d�[��)/U�jv�y1����vF�R�W����E��ƭ䋸!g�K������~�]����+w��G�"o������t� ���ݬ2������C�J0���d�פ�+���B�(vb�p��t�*�zy�n:>����"9s���$��'�L��G�3KPo��j�A��u��Fxŵ伐s3���*S5�^A���!='[]o,fP@�[E�������X�N�#��T�s#�5zYk�]�k�=����I&Qunr�մ�]Í
�􋢀����Q�F9�6v���z}$-��Sl�0��~~.`��꣑о.o��J����������{h��yL�b�:�x+��<z9$��wnݼ-|���U|��n���s8�l�~
��MR ��IMupv�_�)��x�b�j��!&r!\�[I
S+HX���"I�<F�诧'��p��y�$�����q�=��o,��p94�o����~=��2G�$��