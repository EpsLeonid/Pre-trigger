XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C +�R�H�uF�$��l�NVZ��T7O�1�0��&�gs��s��9/����� ��?�jԭz�P�����0J!�tբ�Y�5��~���1�tr����M/)#@)�kbD�'�Ww �e�G!ǽ�oG_u!�|jW���CS`:rrg���fǈ>0������k�ŀ��j�f�A�؃:�U���l��K�v;)]�SU�ԭ*B�v�%}�.��זA}�ؕ6,���wkKBO��%C�KKo��� �^:a��;N�9���b��u��}���v�� �K)�vY�����,��<��+�Y���-
,�o��g�?�sm4�w��s!رfy����ƛW���4�[�FI�SO����� �Q� s7��E��ҿ���)+��E�����GH:
��Ik���~�e�.k[���,�8S��'�|��C޽��`�Rm��P&��n�h<<�)�]d��5����Q+<ksS�/��׏�wv�1�0�L
��A��f4Yb.vĄ*"����ёo^hDw���kɀ��A�u�g-��s��INվ7���y�
�8�"f�a�+k����}�W�fo��.Z}�0�H[.̽O�R�1�B�&B��8!D~��Y:�����b�����/�W�X2���v���\�+Y���Ҳ�5�- *���<�mR���k7�f��^ɮ��a2���a/�G�T�����M�cn�0S�U|��bc.��fVwf`��#p���'��GԦ����P7��V�i�+�`XlxVHYEB    4548    10a0W�V����-l����^��I��}�2Z*�%$�"N�ge�^��Zt��(�o%2 ڟ��,�S�97�CI˖	��;�w��w��2��G�5�lhK	��)�z$�Ud�ׁ��Z��T�x��|I��\rUᾙ�w�k����k�L���#�a"v��2�����5G4\�)��xbO�Y_1B� [-��2�R�Y�k0}RWfG#�t�r�P��u�8H�d���	��!�-w���,)��%�3�C՛)�X���z��yY��U��C�S���q��e�*׿�}���}�����$\�x{���l��"��`ʫ��C�s�P�Ֆ����� �f߼�j:qݒ��]�)M�vh���݃2�lHb�!"����~�WtxRpT�?>|��n���A�ȏ8\߀E,�}���=�F�fk@'zK�^����.����=At��^�i�r�Z��Zo���>���=�ՙG��A;#�3���|�ߌ}���pLg��R��2Ib�o�9jѵYYW�_��Y��宖��O$�\��ӷB���(m�[9��M�x����W��?p��q�ju�L��}�|�z턀+w��Zؾ�3�=jw�)����5��[S��ʒdf'���91۲���IH����z�}�)ܵayA ����N"`�15�~��S4�P�7K�/�f���5�f�f���5��-;I�̃�;����qה�'�`N�i?��VC:�$�XG�5S�hE��U�袧��	L)Қ��H�8d@i��� 6y�\��b���F��[� I f��Y�d��z0�|/����-H� �����SY*Fv�\_����x;���Y��٫���d�im��7����B�9�$��ΟC��5W2dai���|��l{눜��
�SDl�vÌ��y΀�n[囷�F�F0tp��M���M���[Y{7{�|]�O/RJ�=��ocDx���nXa�諬��5vsX�G=�V�"�%X-�Lĝ=�9]�.�a&=��K���-l���Q�S�R��cV�����9O��e?��4J�w���L��?�7��^�ߨк��q{K�� {{~�\]��N�V��\Vh:pR�#�Fx�0]H��y@ҷy��)�^����8*�|�7��>!�.���n�������~�Pfq202�7"��`��|3�"�u�UU��X����>TR��&Ź� �]��
���M�;v;(Ki�
����P�N�3i��%�ٜ���cܯL��］�xg�p!k��\#����ߩG��6�C�h(4�J?�QA�>x��h�������v��F|}�^��T_G=��Œ���h�d>h�ڮ�$NjX����Ǐ`lЍʉFs�cNa,�<�AJ�ҿ��E�(w�u��7		@D��\�:��?�s��!g�x�c�d#�i�>8a��c�^$��H�J���9�W�,����,����v�A����$�w�'�PA+���{���i��gjfx ��G;] z�+��n��gc��H��8�#�����F���;w���|9�s�_e2���m�[���IQ�l�'���[.I��*Pg�f���U�5��uS?��C��Ǵ����ne/l��4�̸C>N��ܮ��6��/��T�.ݜDT^ Q�A�{M�l��C[2gR����V��G���
a�)�+�0��Kx#^q}}V�P���I���X��Jiq4ECс�q���-��*�Q#�@�a���O�k�����@�@�De\��?�&��+�Y_�,4��O%N��c���Z�R��|��Z���0[A�
Ռ���M�����d���9˄�5V���>������\qd6�{sR�@�\RƋ,�5ϫb�:v�f��ǩ��Yw󚖶6�C9��լG��ϻ6�[�5��X6un��Sy���߳�/��7i+���c+��`T!�2����@)[y�k^PZ/�m��?E�h��D�9�3�m0?�A�~m�����V!�3��%�`�p@�	����#��_����5w꾯D�{9n�::�&������4����b�0��]��&lV��Db���z��|��Hdr�\N(�;HlU�ew�2��s��'
}�>�<k�ca2&�E)<IJ����\[�=�M�Q�n�T��&@>�<��J�RߵP|��4Dzܴ���Ng�,�8�N$T��)�ߙ[��$l������ӹӘP��c���(���L���8V�d;�:�G����'�$f���x��O�����	��;�GY3IU@�G�z�����Wݫ�>:���lo֫ϒw��ܴWb�&N�H��� �i��S���|t�k����9�&,�z숓�O��Kd��;{���+���I��{؅�����N}z�G�����6��͵iC[IU��3NA��n�\��$�<=�Л�������!,�G��
���͜0(�*�.����p�\.�bˋS,�e�+nEMD�Bz�2��r����(�����s�zv<���}5���rC������M�(�7�T���S��{;kX��:T�B�ȏ9��-�8�!�q��8����8��>��q~5ün���Di�0v�2�̶���p$g{%�}������A�bF�Hv���bAGƔ �s����(g�/��.<�h���E�b��S�ZE,b�y���#$�W�I�#M��Bt�� �V;\��&������� ���w��%hx��П��Se9��狙'~��X�kRN�	��c�a�Q?���w���	���j�S������0e���?��Pa����3�R����S���/eր�/�~h�-��?z���_~dR��W�gF҆�����OM��"ZCv�H����O\��Rm�y�v�Y�� �3	�$ r=�wZ�l���S�:W�uJT`��^B81�b��S���!�kUtZK�.� -ܯ��� ����^+�}��.�}f~/Q���쐰k��hvb�$J"��)�|���//tg0�|Y�z�&��X�}�;����H�Z@�H��dtRQ|X��	Y�٪��o�}4IOР���#I�>5ǋ>��${�kwŎ�v.�fŰ�������i*�\�P��^	��;� ��חr��R\�̓�J�TRI�ޖ�2�0��	��Z)2���͍����������=Ll�k�T<�)�~� �Ô�k
s�9G�c��D�^�iD�L�^�<b�Q1��sI�=���Ӝ{�� ����&[�7���Bއ�^D��PR:��Ǯ}��̔�co�
~ J>���H�_�b���i��y��M-	�g2>�Ƌ�PlQl��[����<�,�ߩ�Է\K�����7�E��ߧQ�qJ�ٶ/�x�=�.3��\�|d��`?
<?���ݎ�X%1LIx��nv�<�
i�4.�����"�3�bpa�]wR{��yH��H
���
��1�x��Nt�����.#�����51`��\��!=�%&Wr�z+�i�Mْb�����h��u��ï���`H���-k�Np��HLi�
�>8�+7��sJ����������Ǵ�Y�m:��7���)��:ҥ����23��Et9��d�9�.���
�9`�(m��|�tk:��Dk�n�b����5������s��`=��w#�d&�_�� ?��C�,�.��1�e�r�*M2� ���n �&�h�?4;����
�D��2"�H������M�n��X����_��F�B�W��!��M�d��xf
{��$�2��!�8��I'�W׊�% �C��-�|�EP��g�mF�yfQ�+a;�.��aE���[/��e3����'r�'y9�s�x�2�="�Y;��a��a���G�x�\�D�H�Ɵ!�x��	-z�Y�k���&��O�ck��u~�!K�I/��6ׁ3&E뽝y�����B,橜:�$�.d���@o$K�U&��R; �5�zUs�Y��2�@.�d��'^�ؗ�ʻ�\�E����d� �;~��9k����0��ܹ����n@5}Q�!{����g��v�������7Z"�X�y�Va�>u_񞕠]��d��I��҉@��V��^����+v�6��;J���f]
�0�r~�j�ED7|�~Ji���'�2^���E����9� �rs�����Q�n.b��
�x��:�ы5�k�a������u�P�-����y�