XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����.��X�ڴ�{���=Ʈu���GF��y߃�7B�-U{�&��\
=�f<�dcC��B0�/mcȝj�S�qn��g�C�;�m_6PR?�Zˆ��^KkC��J=exH$˛�pY��x���5�;�n&��d�ņ��?I��K]��r%�(�hͽSbَ�q"�̼tM58�@,ae��z�{�ϊ�T&�����t�Jm�F��/��o��6>���|��~f�qW���?U�,�P�,*?�bb=�v2�F���[i�%�8�kzz>9~��(�֎`�o�*��.~�S��Q��mr��JC�1mA}ј�Q�y[��!�n����:5T���D[1�����P�����"����[�:���Vz�\X�`�4U!���`~S����� �NԆEa�^QB��J�iuQHO��,��^y���G�u.M>�΃�:���h'�+A�կ��>�O��߱�Z����EmL�^Fӷ�n��D�>3,;F��#���׻��o��a��h��O_��*��ӊ+��a2�]Vm��'d�-F.���|=eN��:奻Cޛh�Ԍ|I���R*�)�"�0��e��&/Վ������~ͷ��A� ��p��6����M	p����_u��j�J	Q'&��M�@
�i���4W8�O��&_���Gh޻�@Y�.��FU���H�4��k����u�K$�N#��t�ܤ���V4ת<�����)V��z�oy9)D/V.jO��#����I7�x���[%���<XlxVHYEB    1231     7c0��FkfL_�D������s%묐��Yh�����Δ�M2�l2x�#��00L�⌟%�<�k�?+�����Hd��CP�Fs�YxB�L'�rT2�P/�t� �<Ѧ?*U������&�j��:�Zw�jQS
�!w0��i��X�n\�Rs0y��:'���1Bj�v��m���vq^���%"��N۴Y�<��)�}�W㢶�X��X�oS�ݡߣ=dŐ��iF����b�$����H�)��|��rw�{�@�x\W`�jWȁ��B0l��u1�B���&`�U��Y��l%��-4k�����{;]�'ް��㲪�t�۱ɗ�7Y�(y�I��Q~)�
�L����y׉�@�e=<JZ5���5�]�Z��6�eBYDhI��K��n�R�,of?�ju���jlw1��]X���/ꣾ+���5}3���d*f n�L�y0ڔE|п2�Q0G���L��ooa:�����!Է0�D��tf)�8qVo[��9���������>�q�OdL���Q��/y����+L�}|p{���Ơ�G�;�9�b"|�KVW�Vb��)��2��["
�Ӑp��*$PX����b�}d�yX��@O�Ѡbc�]P \�����\�|���/3�y^q�u�s;��Py���	�H6���L@�F��BP��a�.�E�`���|��"m֗́�>j�����	&i�jϥ���l�l)�f��g��/�G[��V�b����]�mF�z6
7<RД�:��+9���q�"4���\�f%���I�[��`��:�ۍ�S�������|��88o;��KL�4�~��I~�7ߢ]47�4]�0N����0������| &#��s��`����d�I�!��������ط���~�d�o���Vs�	�5��4�	�w8LLW�.��f���Iy9k�]��n.{e�Ƒs�Q�$r�D�ȸ�*�q�=�0>f �$Z�Ӿ'r�N��MI�e��r��[�es��T]O��z�89$���~����_Qk1�&�Hd<���������=��(��5ru�PZ�c��M��TGj�/v���[���$�)�!��k|��k�N�����	^J�c�@������@�][;��5�1'B��y�~���#Zҷ?g:&<���Q޼�ݳ����-|ޜ���1�n�Y�~��{�P!P(�wq@\�@���dۣ�k�1islnu� ;	J;��5��B��
���^�Қ��=� �t!X���bekv�8%&``��ޚ��I�tNT�vb W5���r�Q�1�73����5�gn�}�=�\� �^֩�N=�F�a��C�c�,��T����,Đs��UK ��ږ�����>�a�"��n��߱+-���(���u0��'�֒
� �	�_v��O��T�b�>��)���E�@I���UB̧��s_ѽ��W��a(����BYd�I�@�|@w����?�<�X6`�;N���")�Z|���{(̇�&�ȽѶO!������#ꬭ�5�3����8ѭ�0��~�n���U�e�6�q ���N�T�D�חR�+,E�I6� ��`!�G7��&��A��-���HN)&��3[Hq~kZ�oYv0X^1J�^e�"V�]�2|1Q�0$�$�F�è�\�w x3f�둠'�k���l͓�i����A��z���شXԬe~)^Ob�p�!���6�'7%�leHLV��[r�w�����d�3�f_x@\r�D�e��8M��pD##�ķl��T�bHo��'�;i�-l���lS���F�UV��ABʪ�����Ă��uk�c��jI��d6��a��#�~�i�`p�<wHo�E/0pԣ��16�C�p��&"���`�Ɗ@"�{yu�ǹ�Li��G(ǳ9��Wa�-�׆�Oh]�W�\,Q�[p\M)/I0�v�P���s��̶+T%�