library ieee;                                                 
use ieee.std_logic_1164.all;

package Constants is

	constant WORD_WIDTH       : integer := 16;
	constant BYTE_WIDTH       : integer := 8;
	constant USER_WIDTH       : integer := 24;

end constants;

package body constants is
end Constants;