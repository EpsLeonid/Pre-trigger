XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~_"$�,{/S��rLiO<��D�צ�K���UQ>��A� �����m�%Ə�9�7x�g����1�L�J�$������%j?�����e�rF��Īm�7EΈ�� ����O��z��45O脨ş	CUw��aJ~>',Moƴ��{��k���ۈ�t�w�_��FS���x�[�����W�?���7!����j]�k��^ǥ-�z*�������Hv��$�3�G\Ղ�� ���Zx7|����B�R*Wf�FDr� 6��T�g�t:+��*.�2���}�N|�򉣰�e7cCJ�gp��SW%�X|~%v|�W�xsOT��TJ��9g��:�X`3������	��J�Џc�5_��e�11�ء��8x�r����xl��ND~���ͧ�X(�!0�ܼ�L9e�~�G%`�ʩ /��j��˗R��F�'F�1h�Om�m7o���
�A#�Z4gX��FB���id3�1R�'�g�z!��M|�?��hR_��՘�0��u�_��~�,oGɨ���U�e� �wa�I�-��zF|m'#�M�3�/Y�� 7� AH�aDfil5�6!�+:Dn�� ����*��ާC�Y�%�꒪��y�ӂ�N�9M��UY�n�5R��覌nn��6�U7�Ju�|�8H�4	���b���(^i��aBd9~_�-�u��*�x#�����u9�Z��q�z���?yr�)_9#�tB�)�O�DX�<_�u�́��F������6��V�i�����HB1�c�#+k�|���XlxVHYEB    1001     6c0��Z� ���/�I���|�&W�X���0Y����I��X�/NDIc����"���l���a�%�9-N�����|��F��Ǐ=>�^E�R�6��G�r�
?�R\�ט|�Po0���.K!���N%���4C�N<w�9&�4�&��@h�
&�b���#�W�١57�u��3��������v��������\Y�;T�������[�	��C��z�-Z���K�:��	�5ԥ~6]�+���U���5-=6�F ,%��ߕHG����B ,"W���M�-8"%�4���lo�ke���1<Vqp���ѓ�m����if���a]y���Rm*�d���uQ�)H�P�N�>������(�eݳ?���&2ƨD4���D���K�A���J�6b�zt�w��5�jެ�,��۟��[�(,��e0�>�����-$?q�����Zڷ_�w&4A��?��g�g�D�@z�v�����5��/�^9��F��F#��n��4|�2�$,��}3C`F��1�]�z?¦`�fg���>hMD@m8'��m#���8"�ן]зIt��V��,�wܿ5��"&''+�akL�&��^vx9~~�;>y���ydI#��,1�.Ů�E�J�`�=��+8,ٝ�-,_^�tV&_��+����86Q��}?�^:�j%nږ&���.j�3]�ʧ�ֽ��X���ݙ+�U��@SbG�&��N�?\�lɄ��|޵ cd	?�`?��T����hQ�o�ج�d]Z��ә0�G�,��H��P��o��#�0����$�9b����!���E*�z�hם_@9�b@Ӯκ+h�qv�@��xK��캮P�Zx����V�z���!�W@}��1ُ	�_�Y��aT��fs췀���Q�=D�x��Ȋq�_q�M�?s^����kO��#q��y��r�Z�g�q�)�D�[��׈l6|6~�	H�%�Ha\ѹ�rխ��A�R�)�;��>X́�����&����}�B�1x<��1^��y�5:�5�>u�����;׀!���vW��Y��C394)!aP?�j<-�p?'{���{�O]�NG��bv�`���⌨{�,�~9��	��x�����1��(h����I�^HI$s��\���������$; ����Pǂ�i����q<�����o4��l����=1�����#����&�3�le����.�X���i�{QK���}g��3ǘ�w1]��Ki���D���f�3l�T�gaO�T3q�����v.;kY0���1�R��%rW�� wH��[m�K���	>m�n�)�n8�Ƽ�nPw�ܣM�xJQ�7�!� �(*v��5��y[���@�Ӭ�0r�~<��䵼��)�Ș��+�V�z#�f��ȟTȗN���%��6I�Z��ł�*J8�̸�ӱ�Ont�g\�T�2;OJ(�:WL3C����H��+t6f/�R_��O< �^��'������3BWx�g�FV�P8G  ��M�I���tcd�	�C�&φRH�ok��J���’��iǠ�3�,�0J\a����l	��ѫ��zn'�{����� �ir�~��/#�`�|�-8}�U�,a��l��Kh=3母�$�{�|M!F����ͭ��=PV� �3p�{�G�	qF1ģ��X�(��c�}�H��ߤp����[�Ɔ�'*�E�pMw'���څ!6�ϳ�D��