XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���vQ|�f���[郧Ϡ���E��}�{P����Q�����t;���AD4�<��ǩ3�[�K4N�o���A�f�HJL�G]T�?���z}QA�f�C���!�7'\nЅA(�]�5�x�޽sg"�V��/m>�`��2�|d �a��<�6{��I%�P��q�����4>]�$6_����_�f�ߴ~л'P  ?�I����[�����R�.b�ʢ�!�l�I��蔷�{�M�/�2�K�i��|�Y�ƚ�!�NWp��ٹ
	�*���۝+�<fu|�
�@<���
��$ �E���)���f�*Ƕ��J����_L%[9�K]f �䓐��������Iqjz*	�$5��2���$���w��֟@�8�p�8 ��)��}p�@���m�+�H.,���v�m<.9ˤS���>�&�>�\X����I�z�d���@��H�n�k��FQ8`M[���}���O�A�?W�}C��d������ſ��?h@vW]��d�S�{��l��l� ��W��Y�m:;�4<D�P�NSؗ�U<!m��#���sU�j���p
��ѵ�U�#�&z��}#9aLǙ)���c��޼M��H<!��S6]�yo��o��o5qJr��s~m(�52��J�Z���%�/��1��#�pi�'G׸�G%� �Z�xu��*R
Oo]҉C9R�_P%�xd6PV8�逡�4)�b_��M��[�e�G��/n<���Y��N �k��WV��Z�3���ԲF���l>%�e�XlxVHYEB    a19b    1f80�����U�2��C�$��Uc��C8D� 
5ϫ�Ή���w2�{�� ��b-K@eR���kT��AҖ+��nhMk���el.��@�U+��<���
&������X^�����:QE6.F��;�FaҮ�u�7Z�D�x�/�%���K7Fo�K������wg��uuǕSD�QIb��vl�>�$��48��ޚ���h���b�c����̽i!�T{�j'�A��~�Q�#B�uVh�q�(��%���zT�"g�����j戈:��n�d�=���e1���"�����3�e[�8O���c$*'?�����˘3���HM�+NGd$yxj��:���F��1�vk�ͫy�Ȕ̥ȅr��T�S�[�NXS�����T��\��x�I_\�����Ȅ�%���1f.���X�Š�EV]�yY�������.��.l��;Ghڶ���������}�=��o9���H9Cy��*�<�5@�%�6&D�d�PM�x��)"���G��}��׌&g�F�/\D�z��9p7��ģ�`e�<�++0�b:1����~�����=1u�8L����}Ď�
a&U�R|�@�se,&Z��Ed�X]ՠ%��>�,��ȪW#H�
��A0Lh3�:Ƀ�����b��6��������[�ϟ��p.~�q�H�*��Ѡ�{��s���ԧ��8����r�31��R{���5G6�gV>]%��.A�ҏ7�܂	��N^��4f��~�<��]��$��1�c�<��O�o���^��M ��Z̥�&(����zLr�Su��zTJ�aT1M�-ˋ�9�e�yXU��d؅k�@���ه����������~���Ӗ�<[pf�����(�Q�Hf(�W���ŗ�������گ�0��R���n���z6s��,����m���v՘ʗH��gs n"RGJ��DYk�(Xa,��������a��(�.u�\2Lp�z��3C�{"l�Rs�K��KPD�eM'�c=�57+�q4�cXo���^߹���9�wI�K�u���5<����(�C=a��B������b�G�Z�L����a�Bu�;�3�p��[����Prqe�X���/�aHN�l��A����BΗ?[~�8
�0;��@�tGj���
AA�K��J��w&p���S�� R'��c�&� ���MB�aI��-���p�\�pq��tZ
�O�c�[%}�1�#%��oǘ	C���� �&jC����	�x����żc<?Ҭ�UŉLL��_
��K����8[�9pᤒ>=6��h��S�S�@>��w��r�'@�,�`�Ϩ�0-�ev����QP;�y�~�@w'I2��ƹp�b��(k�P�=�[�K	<�v���9$�aQ�����{(�JcS��ti����B��^�ܲc{����e@��� -�MLw �٤�7��$5���M��ۥB��[��#��uM� �����7O.�ǖJ�6sHC����%Aؗ��`x��u	q��V/�!v�Fy&kċ��AGVܭ7�@��_�
j�����樺�C�{?��*��G�x���b�-˔8K#�%�E1�:�>�ȲCs��g��ה��+a�-S�m<�T ��]�l�~b����O�l�k�]#e�W��K��.9kG�����|���f5��3�\����Gx'�~9���:~D�Tn\TD�D|��^�G����:��i� �+,����4��k�|��##�i9�ȟٰ�P��KF����pR0tL����GbD�D �`�u.�4��>4�kj�^�AZz��@�k��]w#��s	=� )�A��b�d���S���_��!������9U��r$
�ޔwdƽ;r���s��Thluu��$+��z��ޫ��;R��J �ߋ���_a�ӟ�8��"ӊ4���җ�_�o�fH/wzd�!%7I��Y�~ cA�z��}ƌi���=����e�6����eN��#-��G��T|�|�K_Ӯ���� A�i,p����`~������5�τ9��4~�N��9������ q7tSV��tz�Is�萆�L������`3����R����l�maS�R�/H��Σ�5�ډ���!�nlr�[���U�e����#y�4B,�\�l��A��B�������"���~�3�/���T�Bs�B iW�� 
�#J�8�������'�?_`m�Έ�4�B�!��� �@0�����b��Nq�avtk�ɬ!��D��H�U7�=$�~=�=�L��8W��a�U	~f[C8ƨ޹�����qz(�g���ٱ��Xf���'��v�Df������e85��o���Y�s�&��n�>|�;��B]��w���5@�Æ�lT%�x�������rP�y˝������HdF��o]�#Y�����'�4w������6w� ��'?��J"���Į�=�|e!����1*�ҮF1�qlc-�:Q�Z�3
��0����ɩ��R�7`;M����vz��+��4ih�8�8��U~\<���Dv��^g�ٟ ��{����_��ھ�ܚ��i��\�<c�Ҕ���4�f�i,m*!@T
S��G����2<�w���t�dҼa���go�ո	Yy��;��� ԛjWh�����囉\��=�ۿs�����g����s�u@�EY����SїRq%�b�}�Ug�i��%��]dp��Ah�$��()�`������m�m�S�8�0	>�պ}IYﶄ�gX�NS���7�Q����Է�
]�8-��
B��!�dpl����N��$��p�$�N@�k�<~��#�睹2��q���n,a��� !brA�N��(6�;L��=k��ܖ��G�F{�E�Y����3z���1J�oRݦI*�v���TP�R.��wl��"V�DSX:��4'2Q��Oe�Cyd�Z���7)�:n�ď� ����t�[:E��{S��yWs�euѧ&"�X�~�;?l��a�s!u�G��HP�c3X�t9����*ɳzԡ��ٷ�
;�^�.��������e��<]����߯�Ch���dJ��p�%���DF���2� ��
ܦ�;��F���4�^���Ta��$E$@�C��E�(����b�w#K�ű����(;HdF,WI�i@eTE���j�����@Fm��a��NTxbzX�VB <"�m�k]9�YJ$�$��W(um�&��:yS��P��8���"w��qks;Z0D��C��5�\�BY��r�%�`���Rj;�s�o ���H�/�_�d��[�e�8~lʳ(�/
�%��)��b�x,S&gV��SӐO�b��i� ��^ha��b���^6�s���܊�P��+<VÝ�%T�YJ<���9��u��Uu�����D �P�F�����sb]�p�/��!~��)�󗕴!�5�>���~�t"t��4,$�Т���h�/�m�В��{ Y�H�<9S ^y���vVCHca�n}9�!�,T0RYc�*�Q�ZDM��$�0�P�����I�.b� /}���",�oҒ��w���l��K�� V�o�?B�M��눂���P�d=�x�ۀ�� ��0ta�_�Z�MSqm��N��������I��ɕo(]��3a)�G	W�O���^ߦ̘��Q~ XB�:�H��!�S���zF�[��N{���-eC#�����(���]���#��j:�*|z�i,��'�����@��Bv�ba����Aaw��FD{�:6�D�V�llu��S#��NJd<Vڋ_0Tߺ�vz"7���1��V��e�#Rw��p�)Y.7�ؼc���J�NGa��8SYkw�ԮV�%����Os�S����RK�h�W��'fps�K<�������!b�6�c���ma㥼|h(�e,]�'�}�����:k��z����u�[��ך��Dz2fo��8�XF4G~qv^A�bPc�l�����<Rҍ��ʮ�R۫�Иx<شDk`�Rkb������}�҈z�g��Z���?ī���\% Ch�@߸m�ԑ:��n"h�4㯢@S^Z�>g��SH.w\c2c.�Q�t�H�[��e�K�/��Hc4	���"��W����V����ХLq���?f�G^uW��^�YG�twZ�!����YI<kr���
a�X�f�� ��I�1q��킛�Rr�:�N
�	 P�����-�.�z�V.� ����-�w|[����5ƽ��4P�[�8t�#t�6�Dpl�WURg�I���2�&� +X'O�TV���Ӣ���4N� p�n)�����麇C�[8�l��Bb���qa;�����|'��Y���m�*��#۞کI�~<6���d�ݫTY>� �=O;���A��n�K�I�(4-K��}�Ӭy�ǹyGo�(J�E�)�YSU��-��*�ˇ��s!�;w���\��e&��F�&�538��fge](e#��OZ�֖0���s�z�
��;�{I��$l�C��N�"4Q8��5�\D��Y7hFzi�#��I���r>N��3h�O�$h��7��@�ي�>��ܮϔ�nE��'�NT��T��܂&�)���m9=w�c�uAyp(�3�叵I	�_tѽ/&��67_h���QP���(g!�r{�|!��O~�1����Ă���� �Ĕ�v�d Ʒ&���_4s(X��\a�|��7����7�հJ��c��I:��[H�M�g(����?����[� lY�z;�=UHK��N�s�	�w�)0I�f���i,7�*g����_�2�HW_'ؕ�e/��O:''�!>�+ƝU���&ޖ��j׼�w�mCh�a�����G��녒D�,�J�Ɯi�k�������eb�š��	�=��"0�p�5@Y*"ѿ�Q�9�rq��=��)�}F}	���ċ4+��rV����{�SC�Sl��y��'�5����_������_+?�� �ֿ^����d���Hi�W򈯑7���~H66��*�����$�G�?� V���ҚI���-�M��ѽ�6��m
�܏5�(b����h�ی��'����e䐜�@�S���Sn��	��@����E�w��5Z��_)���LX��]�m��}�����f3>f����]��bp�KA(l9)��[Or+���.�<��Xd���.����r%�Ap�d2��m9�Wv��dm=`t0�5���0%�^"��T]���D]^/��Ҋo]��F8�B���O���tG!y��_J�.�G��� $Y��%`x�oa���2G��__7��7��#t�X����F�ꋲ�vyb���)cH���-��j4�ԏtE��ڕ��P�;�#/l���ҬZ��.�V�-�2�ʿ���y㪒�]b��@]`�1����6�-��a�l�z��@�m2�`U�NA�u��+�?��n�����M�Pi�ol�]��9��͒#-XƷ$�����K�65h�Lu��%K�v�C�<؅�1��j2߶���T�����cwWH�#�宅W+g��G�6��7Ғ���)܌[�q�n<���!c�y�;'�k��p^[T�2lFD���ks�����c��Z���U�T#�&�0�aE�8�% �C�}W�Qk,~a���Eޗ�&���`�ț�	B_�<*%�#��EK"�Ͼy�h�,������-��%@-�����G��d�=�]�l(���(�_[/T��k_�Av�*�T x	L�uVI�+����@���Hu�E���
 zn%�^*����b� �pz�⏘�t�{��/�^��ۜ�AŢ,r�W*�އ*wb㎝�R�ט�h��s}�:������𨇻�S@co����������D
3J�.�Q�Y�4�F�\������X{ȿ���XV�C��n(�� )uK��Im`ω�|��c�-������پd� �ե��`�:����������2�HV�����|c����x�^\�F��옄�����.R=cA�5��ȃ�~
���������qYS�3����ݒsOr������i\��V�b.�v�Qߗ���hf��Q֪zx'$_/��c*Q�L�x�b
��E��4H�~%��N��F��F(Ot��A��3w��,�Է&f���"C�Zd�P�z��Y���y���eW>jL���Q7�u�r�x����B�b�q����Fwg
+M~�5㫙���3Is�*�*7iG?��BSҨ_�ߝ9�jl�4���D� �5��W��T�u��S��{7HXu3gKc,{���Re���0@�`��Q�PNt��K������*7x���5 �C�n4��3��T�����&�>\����]�,�Ot5���k8÷	�E�#g@A-�Iυ��)�J�-.Y��1lɲ��]I��RW6�"}��u����X>I�1f�i�"P���R�����28v���P�7/�����X�p<�Ψ�<�K����!���&_Qi����y���9B��*9ĽmU��lD���Y�HKO{t��P��`x��� �+g�����	��CT醒��'�k���X�dR��j�@7>�ē>����Lj����	�Z�Rq^A��8lF���D�~9��ӆ�����^j��He7] ��@ ƶ�*�٬A��`�Һw�s�3��VE��Q�����z��^��
�x����1T2�,E��?x�����y.L��U[���0����!R�� PC���zD��c��D'9���؎�T�&����ͩ��I-��2$3vL?)��C4�F�����t@{�x���WJ[��Fym���V������ο����j��29<R��9HE�{{�A)��'n*[&��IJ^��`;BQ�LLRA����n��+�B`xs�.�3!�an2��<���~���:�ҩ�"�d?z������{� S�n�dW��' +V�U7q�MRvs�0���9�q��!p���A����FOM!�Z~ ��}�>�)!@HO}Bu����x3�{H)�M�Y>*G1)�,\������������"ctv1,l*8?�v�����=�+/��i�@���U�C������C�d�ƻ_�O�4�V�XD�q���[�[����;͹�Ec۝�;�zm���Y��g� Hj��Ń�ܼ�������&���YR�ƕx���M�D��w4}�˯^w],�@���lv�{��}��p Y�4�\��fV�Ch鎗�Ԓ����&CQ�0YAAABɌT>ZP��I9�v��EF�M4�>J�9��=V*Z
�x��"�u8��ڙ���~kʏ��n���;��u�l�Ӊo�������K���k�SV�.��]Ӄ�f&� c߫��ok�Y��{�>�uR�g>�EJxX�k�Cˆ�DM��)8M-���޿���Vg���@���fBϔ��a�D�M�(�m���&�a�ݱ���H|��f��ڋ�+z+}���ۇdr2r���#��=%W)ѯз�|!�M;��e���f�ϟ��c���^wIZ���AW@`%�[�gzK�+K���î�^�|1�����jO�~�Kg�J�����:�##�F��L�&Y!x�L;��l���,3��,�����8�\>*�ы�n�� �'=YP�CGެa��$�.�lʢ]�U�����r��������'����uye�>h�D��|��
���SC�A �y��&ݒ[��'気=��28��Jsb;����������a�D���c"2%�!���F4�u� 6���g|$��+�||Ee�d/��e�om铄+r/Q��k-;��܆�i/eJ�LJ;DQةy�QT
3v���0�UT�]�Kp���E��ka[E�f%kufOT��K������W�D�u(����>��)�R�Z[~��A���*�36�$��^?�