XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������M����s;d�ꕤ~��X���q��x<�d��kx�,I��jɩws
�,Ku�1fZ_Ȕ�S��>� ]*;�1y� �#{y������L���HƋ�i7g�M�s��d�x~����2�)��5��x�f��UO��%R��|�w�h�h�w>��������CH�b�V$
:eePX���7/l�E$&�%q� �N�{����i�6Qu������}����a��į�ॺ��)�,�s��۔���`M7�;ăo`�����~N�0�r2�����/��>���c�J�7��x�r&�7w��K5�О���M+�J'Ԏ����tL��		{���#�M���!�d�9l��Q�He�_�c�i��s���eDnb�]����(F�	�T�ka�5+���bWr��r��f���\�Ax,�6� ����Ls���pȟ{��|o��	�\]׺T,k�������$�:Cq�9T���[������q��n���åIGӗ���G���fv�ȨZ0*Y6�[�����)�Y�Pup�qX�3�˓��F���`�_6�7��c�c%�G�,"���]�����[ӓ��Jӕ��B(zϽ�m�K�~�.���5QJ�n�3i�,�,]�SG�Ȭ(����|���T�A�_���4c�t�ꗋ�h����an�Ԣ��eL�.I�2����5@૟b�z�h��Sl�c�杉fV��khȯ�s���LH,�nk�ME�c�:�����XlxVHYEB    523b    1130�Jb1}��C&8��"6ᕧ7�>��l�?X��y��ӭm���1º��[
���Md�1���5suv��d��ph�N����J�3��m�Yx�2�p9��j��F��Xț┈��5�K��� ȷw,�E���F�]Kb�n�]��Zn(oѐ��C釴9�=X�}j��S��0N8�"��(�tɵ6cЫ	 �Z�)��_���moъ�`��ד���l���hV��ԌK,1&SYC��6|�'u(~CvRĮ��%�[�.�V�X.3K�ѹ�f7n�qK�ZD|��cu�`�6+;��cY��
�c�*׹�a��x5���`Rz����i��S�,)�����'���_���!�v�AU��R%�:b�a�19Zg׸�i�ص��,&^~�gEe+X�>��Q�9��$��*����eD�7���T��I<q�	&ٰk��4Ţ���o��F�eJ���@s��8٭T�� 'pX��:�����z�Mv<4;|]-��6�$+��bV�\J���b���|���^�D�����6y��o��
�!RPs3Z�@�2Y��4�v�M^|Ffژ��$�hI}�VD}6~B��/��17�m��=(�q��f�F���P:�L�Lc�������ɦ��0�6|@�2q!k��"|K�:_fwE"��i��͏����'dF,jG���yF���P�JcK�=m���s���l_r`!&%���n?e�#��ǝ����Ja�	�?⟤��.u|�N�K�=�P�.9U%�C�Ǌw�Q '�Co6��n��o�%1R�D�g��O`|��5~�7ӭul�2�61?9��#,��0�N�|��:�O��|F`1���WH���rHY����EGv�B}o�7�F��:��(��6>������1�y_QH�Lm���5O�O�WVbTG�q7K�mfc�RO�T+�����kIH߿U~�j�-͖��~���=8�RbY����x�z�(U�+t��������/a6��c|>5?�<�L�l�P�7��l�u|��:a�/d��m�?ͅ�P�������1"������q��|�D��Q�2r�eje�lWN?�A�Ȫ��<�4�y@H8�Q0ч��� �g.�Ɉ/��z6��+fF_Gͨ��?��2�d��+��Q��L�͹���ˉ؋a9�>��+����]"�l���\�6/����m�\͹@ �5�W IG�3��P�u9����%�4V:��p�����%�U���)�nwC��e�k�!����qY���pϥ�r��&�A��zd�j�0�z�u���lҾv��+f�u�a4��M��9�:\�ഀx�%�`�8��e�ݡ@��\�r1�@� K�*H*-�\-��ý���r0���\��ضX�@T�RT:�и����ê?��\t#zLOy#M�K�;�}��A눳�*�~�Q�����և�K �(; O��E2y��\���ߨ���󋤢�TY`�4&
o%ai���_Ͱf���GL��0I��ZҺ��0���^��@n�&��J�7&�EGzWݙ.[��	����ݩ����h��4�?��ir���V�啝K������~6�w�K��.���1�]�_Q=Q���Yɥ.��\�q{L຺�PV�__�qq�&2���Ĝ�%`o�KV���������Y�Tģ����n�B*iG��WXs�P��v����r�ze`Y�C��JvQM-�(��xU[O��G��D�=��=�G�~�&os�ۂ4�a0i���p>��Vv̠�rx�i�"	�I3�����Gt�G�Q3�A-B��_�0[)����	��71��϶^7!Ts��4�z�g�$� �l��n�Y�-;�K2J���1���rϖ��4��F��
q�- ��3I�:"���pS2QR�!j�S�Y��`˒sݔ?���b����X΄��R�H�Z
r_(��bn�(���Z�i���d�H�xL�W��5�n������}�s�͵�峘(��T�5ڱS�t3����^�6Z�IV�#N{y���\�-��k%��(�I���osN<��{\��S�������H��@�t�Ƀ�YE�w��a�1�x_�lyVq�D�o�p����a�Zʆ��%3d�}X5�h�8�"��o���L�~��>�D�L���Z%=+p2�Y��S�1�� \���{�r\X��>�A֚.m3~in���6�u7w�\�������Ԛ��9���c�^�g���o�L����ł�G�h��,�1�����\$��NX8/!��}�9��J1ؖ�n�n4/��gTձK�`�1`��}�5Z4p���tĽ�,��!�2���͍��N/{�zC�.#��XI��1�l�H���]Z�,������3[�n�^�i̙d�肉c	P�r >�"��I*<� Tf�5�}�[�4O�xͪ6�C|�j �?�Z�9X}�[���@�ڧ�O�N�U�S�����ҽ�.$�N~�O1����LW�Ŵ�z�\f��3�T�r�����#�/Gb��4��v���l��˲�ATl*ZN���D����>�*ã�C�ł�7��1<�E���b�@R����}1(@�ꅙ䮂.�]�?q��씮o$�3<5���*���ď�j7�K��v��*�j�Ft(�Fk:`�.����Ci�����p���jRݬ��.������Sz7��>���?�e�,J�w����C���{�`����@zwHpW�����O�n�O%t����Q�RLp��ԯ];�6uO�I(1�2�
Y*�,����R+l���s��C��H֔<�K�������,�)���g���S����;�*�q0���Z�����f�v%�q��ڪ�w�8(��U���lRa��M�bA�4�@P���52�o~���j\22S(�|�x�&݅���U��ո�ݹJQv:Vl��U��>�4��09�����r��^���uP�xB)]��Z(Mb+t���*�D���J�s��5u
u�a.�)����͝�J��Ҽ��Gj�M�	2W�a��-¨�G$��t`n�.6�� !�˟���=D�DS��kb'�k}��⨫f���+Qx�	MJ��v{غ�"*��lɥ�U�L��(�����&*�Q
��a�c�n�����6�}K`$���:��J![H��'?M$�̲�<�Jmy�
�芓��K���额4���5��t~5y�T�@��d9�X�Z��C�N�߼�`kF�i�cӆz�k��M�t�:�I��G��4�ld8�]�TV�l�Ď��z�^g��XK%�u�\���$�#` x�LX���:�R܉�����W���L�X�wE���V]�#c�
�\���¨�v��fC�L;���z��w�W]�$�d`%�!k�t=�Q��
6�g%�����2-@��^��w-|��8BYz�u���]t�!�mL��������4��jN|�S@���U����S�t.�\M�=
P�!KN�FB�ä��k��P�l�\晜и3R\����822�֭�D5��1U�WUp�+I�>����B\PEO�Hp��t،"�}ಫW�������VB�Z������)�p�R�
p��
c������YF�_)�m�h>�q� a��	Ud+�����o��i�t�x�\��-�e�Ƭv� A���/j���l8$�{�Z�Ƴ9��Ј�+�_�
�ع�������&�鏻2h��v򩡙lЍ7��J��$�ڹ����2��r�k;6t�v�#���ק�-��������٢�����E��<5�W�,����O$_3��%��*q�"��Bف�J����%g�����rR�O5��/:�%�JR	�ү���&-�5�!3}�"��}@RXn�@������gw�fp�W�������T�V������݈��Я��)}�%���n�\��E��̨�/FT�ҭ�F��6��(��{�!ח���qv��X�3+\���Cױ�1oB+����3�6�%2k#=ݚ�����TB��Q�8�[�x������{�K�RƢ���	�x���\����'ʐ/o�\n����(NG��(u�쐇��L�L�r��&�a�7y�����'��JMa͆��|�-r��i�!�@�4�V�o����]�N$�}�Ti�l�v)|<��WH��`2��e��.I��Ks��~� ־V�x~P�S՚A��,;~�D�뭌�N#�'����(�D+��Y�=U��;���e)���ӹ��[�A��.\n����t)�Gsx)��=�#��i�r����w�7z9O0�&���y[+S���RY�LO��w��IB����[w!��8jX��{��R�IY��