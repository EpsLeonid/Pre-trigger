XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����|;ݣ�����>w�yGXp��f#�r֏�)c"np�D����hg}q$�r|,�wr�#y�����hm'8I�!iy}��%��IɊ�x�w������2���B��gwz^�������4�j�u,Z����N��%l�s�r�<YX?�DL���>�������J�-���5y���p�C�5(�%��(a+f�4��a�X2�d���r&~��F�4\�x��Px���_T�}�!�H4�#P��;6���4��2�f�S���^��D��ͪ䩜l�)> I��]��}�5�x$꿈���p�S?cu��k��ñH!�qEǀ�f)y1AN�s�������&5AZa��K�m������I��YGU㽀%E7_������8�fZ�S�}]��lz�:�4Ȣ��`�0d�.Q��4+��)(�����S����cLq�ˤQ�M�x2��#Z��F�3�f].����n�I���3[���.��0�1��Z���b�����Ú�[=�sr��Y-T��:X9\�d˭җ�����I=��Z�F]��do�A=����S��֑��%X"ֶ0Xٷ�S@�������7tԔ���f+o[�m���΀�,٪Z�B�D�,�W �qa�3��p��3r6��X��T� �m��x���?�~?:�y���<b�f��1$�� ���ݬ����rM+ѷ9���C��m]�`���Q��¹��ͅ>w��48oґ���PRy�m=��XlxVHYEB    1d01     a20�♖}�2��٠y�V�sZAC6�,E��	i'r⌲Z�4�(|����b�U� (g������-��>��xGJ��%�>1���¬E8�t��;��1S�{����ˆ�/�I�v"ܧ��`'
���P�&�ߜ��Id2���b�4�g��" =q,���������Ī��ԉ���AΧ_���]��N�ƫj������T��H�%م<2d���7���W��9ú(--bx|b?(���R�y-Q�P�+��.5�c]u����B^�c).D�G��58`>KԴO �@���s�Ԛv>o��@�����+ŚX�J��׋��,񙇥$�j���y��b�,��"��B,Z���6�.)�[L���V�hٹ������x=�&@Ou<1���[Xѿvuz���#3�0Ґ'}���ʝ�r�إ*�3EE�j y[g]��e���{H͍P[CKO�ym/�Z	��ϛ�|�h��y�K��s$><ߔUq�m�79�.�P�qv;�Mv���v�T5[����\4�N��=� �l%:_�&��D�����.�N�$�ax��\7f�l^���<����sU�3�����U2���imI��M],%�����n�g��g��}���0/qb*͛�2U� E�W�iI�c�1y�g�f�^L�2�Cǔ26����bDih�H'�	��\�҃�����@��f�=�RJ�̀����ߌ�t���7��D���1�`|�<���}h6\����&JԒ��TrU���X�4����E~/�U= ��(j�(�%��5T���v���Z��U
��J�|�k��')KnCB�`��̫s>���%�C�'M��]A� �p�z[a�uw�ݰ�z0>��r�����e��bF��t�i��UՏ� �T(�ĝ��kT�kl�2�캱�*L��@�	����b�N=���-H^�`�a1RF���",�G�&�N%��g1�Yn�5K7�4�AKxB�f��d_���-K��:tL,���۰�Y����"7��ܤy������	',�~�u�.<�zI�`u�Z���|GQ��ٷ��ޭ>�w��@�F<R+���]>�?��	�+����YR;��Z^�i��֐�䀉1?֮h��,O�њkC�m��:e�T�Y�C��|��f��8��R�k�8.gD�Y�qf1���#+f�I��=ż�a��=�GL��4xD�3��½� �:�2�%ֳ,��\�e���a�|+�}�f�0�26IA����ǐV`��e��>� E����^����T���Hs�X\�,t%�ݖ��g9�o����XfJ�]W�ߖ /J[�}��+��vHwS�;1?��m�$<��U�d���<KRW��&��,J��
*7��4�\��O_\�״),yC�s�=e0���k�4Z#�V��µ:<��#K�q&nƥլ���d��ǌui���S��T^5͇L���C[!�D���l@ꆩ���2��@�M�(nE��Ans����Υ��R9:y_�1I�0��� A�B1�e�˩����B��ɦ��};�w�;G�| �\~������j����e3@�3:s���l(�3
�Dmܐ9ڽMrA$R9����q\���Y�L��pٺ��r,�gS=�5!0�B����Y1����q��%�lG��n��N-Yƴ�((��LC8��/EHRv_@#`؁�/�ßr=]���/k.ž�̗�m|��G!�X(���O�p�}}�R�~f*��	rz8wx�wʙ�k�S�Ɩ|��}.E��Ss����
}{.�]��,6��3�1j�Y6�3Oh�q����g}H����*S���ȷ���(�6S,�o˩Hc�p�67&��j� $��m�lѨj{>�8�}/S������`���5��l����D�CX��﷗ �ԇs/hE����U�}*F>lz7**���)�V�Qվ���W�W}��=���;�Dᅆ�e�o��Z�E�%h�Z{ �-�����X���媨;%������M��_����{��eK�a�Z����ɫ��$�e�	ژ�cKk>�(P|� }Z���Qdo
�j��n751�����&�ݞ�m����_�sF��8TZ�%x�*���#բ�H��N$�]��W��9܅�K�Ld"��>��Q�nR�����J��,��`��@�� ے&"G�������݋��k?~���K��R
��m��2S�<T>��}v��ִBiZx0��!�D����>�n��3�Ԡ�ʥ��m��7�I��=�b|�N��d�dr���f�E^�3��X����!�=.��Lv�L>�2��v.y%�~�&�1Е���7�R)F�X����>"�da��v,8��\�.�s]����׋�up%%B$�� �O^�j�3�߅0i����������J30��S�J�LY���<'�LA�65f��hY�}�{�_{�&"�8����x<G��u	����A%{!�2�#3g��?Ԟ�[ia�_~y�N�&��]�s�ʨ����pp�s���Y}�N��8���g���