XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���h�4\��Fc�?�,Kv�G:2��/�`�;�f8��Da(I��ЇY!G����DMq��*Sz9GV���8�z^����yG�4ܯ�V
����|�t#���PZ���4y��|��nwx����rgg��n����QE�@Vߞ�|�֓�.u�o~�����͚ ^�0
>)�ʘ�ؚ��u���{���ޢn��E/!��XNDF���ք�GZh�3�fA�9���)� 
��E񲠌�k�F� ���71+3Y\�
���`���Ơw���P>���8��&�D[��禖��u��ɣ�f�~��B�47�yȉ�VYY�V��F����]����N��@�#*�|�POc��k,$n��/���U�����(��!����;u���]��;�S���wF�Z�8V Sw�}墲"cl��_�A�y��q�C#�k�Q�?�2�4�7��R��&�7�+E5���^�vw�2	F<���W��u36��iT�D��[s���,��\�����/F��EXb��Mt3��܊��4�b�I�Zְ��ꄋ&L���IY�Q�e���`��d/,�����W�Ȼ��O��ra�>�n��C���E��^�_�P�XK^(ו�A`/�����1���C���u�0|9T�]b?Ie!%)^���`�ySy����y9;�}4��R�}Z(�W��1���J�u�"$�?����Y+��xϩ���FZ�I�	�֝�.ڟ=�W[y��<c�*�t�ܥ�~�&P�]߷�j6�0XlxVHYEB    1017     680���H�cE�V,��r�V%���
p@H�IA�6~e�;x��x�ף�5$�f�b����,�r�Q�	NS=�Q��f'9�����+^k��?%[Y��:��o�����`J��&t�qK�� ��?Ͷ�8Ur�ܱ�'n}�X���-��+���K������NqUx������P�7+��^�
��B�OQm�M�Ơb��N�u0m t��x�eV�w�H�ɵ����8]X[��S��B�cq�C5�C1�t`�'����4�]n�Gx���\�ǹ��Cm����i�n�eV�tt:"a$c0����[�`�ߌ*�}�J��	3�l5�]�2@h����t
���8�y�R$��Ђ�?�C��(LpF>��Qm7V�0�ޖ�!�'!J>	ֳ���h��DT��`��4*�J��F
�&���P��k˻��4PFv[�}^f�_�筐Q�2J����O�"�0���O��ۓ�YÏ�����>���io�����J���JL^A>2�ZǢ]wב=�dY����A�T8'�4���ᐮGX�!�Ef�}p1���}�<�'����P2�+��S3U�T���k���AT�����`8D�G//��j��-���C�����ru|�ÿ����:y �[6hmN>!Fy���NF���f��)��QFC��$��7��ތ�S�}�xb �=�~3G�>�ŻH��[�x�t��M���T
^��H�WYy)��$K]ਫ�Ӣ������6ƴ���#�F��m�0�k�-�A���IUٽDA9e��ݮ�JiFP���՝��[�x��yo#&^Uz]t�+�9�����"��J�X��T�;a��;,d��$tw�,��� F=�z\S>��0���� �g�l2����#? ����Q]�cn]�Rҡ.���#�FK�� tcn+��oK�3]��J1V}i�~��2��ߛ�E�!�YO%������gn�x( {F��X��K�������s6�N�����0��A��ћ��nbehy�f3�s�8�5c����Bv	��d	�{��DhS��`%�C�(=�U�+���K7�� ƀ�@���!u,U��g����+�����E^�� ����Z:>X�{j�a����җ��Mdh�dhJ��-O��)�����G-� Z��.V�?5�	�K�k�>+�ͨvD�I�Md2��ׂ�cy�	���ͽ��6��}]���T�)Z`p��|���x7T\	a�����Y��!.�
Kl�9 ��Z��x6�T�.e�*[���6�>4jg �F���'f+�{�)�R�ёII��i�r3[�@m�w�u�E&�/�#� L?��&�)�sʫ��ډ�q��g��B���)�b_�JUB����1B����ƱZ��f	����F ���J��{$��ۉ`�s4�~2���Mli*���Fk�A�Hq�y#�/r�NA�� ��,,j��|�)��[���Yјʿ�(��y�8'�����(k
��"��Q�]*3M^����%P[C�H�Lۂ�LW�*$-Z�5�Q@M�~Z�i��zB "�[A�����]F�/�H�u@�V���2ls;>�F	� V+OkmP�U��	�Z7U�͎�q\���w
���D���"cY�䓢e>#�{���+