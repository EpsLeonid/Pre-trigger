XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��n�~�R&�_�G��нC�#|���L��jEl���0�����FFU��������:};gU׍�*��8(��ݲ�dd=q^��t�9��s�Ulg�3Pp���в:Yݪ�s��@*��/u9���ӟ�-�aȞi�d�F���'���Y"�a���-D�rkj�u�ؒ�O�ז���l)�JK,E��Ve�S1:��H��F#�_;��"A8�%�y�v����r?K�q� wr%�d����[[���Zz1����<G��\�uAhv�Ѩ#�^�IM����X������
jw��Z��fO���o�i�p�k�FUt�(K�7��>�n��eNTi�+�4w�?�p4?�|�5�V���&�8��^��f?��!0_|_�?���;,0�B��;����A�F���ON���pe]��W<����v�9b>�/p ��J����C���Ğ�ΈC]���{��qV
@b�;��I�m�9���� �#�T����|�feܳ���:�	d���>�p!�^�����֋���6� �
��?��������t>��4f�~xE��"aM$�AF�E��_�P̖��{�/���Z�K(T*w�8�����_�nY����%��L|� ٱm�!uy��g�jL�&��P���9��쒞�qrD��Ƽ}�1!�g�Ϲ}影�n��|�ɲ��P/��87t}3ܢ���w�59�`�ŧ�����^��b�]r���V��f"��j��dY��k)O�U~��XlxVHYEB    523b    1130`y������o���Jl�Ef�6���_?B���j}i"��A�B��!�?���dJ}�u���ZtP��൅ �L�������K�;]��ҹ�AMw9�֭I��dOcc���j���1� 6�E6?�z�ـ�%�$��

��U&��s
�8_�Z_$VP�nE� �y���ǋ���ܶs�Q̍~����V�JbK�R�{J�}A�Wp������6�S�z��G���"iN��k��l�Wq�w7�9�܇Y��ղ	��lcC�荒��PB{�o&IqF�����D���<;��0��l��O\�����wl`���D�7�[}�ncS��O]�����x�u��eU��/�ז��ҷ[ja�7֖�����qF��ѩ��h)Em�fm�i>BDuڗ� = ^�i͓��Y�-
tY�&����tW9�1n�s�2k�g���e�<2�k�w=E�m^�I��jYˡ�yA�?S����y����0C,��XÒ���B��ӽ�2}��%�؄�\��|y���d<�^�_��؊ԡ��>7�C��2z%��S�2Ϟ˄p>�Nz���PK�Ք4���F9���ʛ^1z�-Ԏ\�bj���3��~�dO��{7�`k
���b0��e�lR��)D�ެ�O�f���0=V�Ŀ�*�SL6�i�O/I/�'���5/���gf���P��]�����Z�J�n B.����}�}����S�JQ�Z�s�<�����	��S�^��@�ɃU���mh�^�|c������<�G�.[��R�\�`o$� ��lq�/fD�ʘ��Ku�1\������n��i$%���h�jlpl۾��}h*?/�=�V�6`#�P��Lx�F>���ȟ�~�) =>�e`���_��\��o��]�e�d1*B���<���AǸ9��s�Ս��.���θQ�2�DͱY"�c���̰�����i��D	�>1L�Dk.�����Y�TD�t�z5"����x�,�J&AÜ���������ܭI�>tG�2
��F~��ް"}ۖS����D�Y�)���`F � ����ߐĥW YJ �@��5����*j&��P%��b��u�ϼ%D$l�q\����6jx80n�N�� ����F�e��;������Z��b�ӫw h��w�K.�����$�u߮�7�`^��C����rz���vF�� [�XmD�?;���椴�l�۽Go�aM�ɠ$j��ekD������o�e<� �#����-����֋���+��v���H��ws��kӗZ�����ދҩVǿe��4t����}��h���w��8-�h���괛s���$�bݎ��=�_���n�y�����,�X�@CeJ�(�^���+|S:�04:z���oc�����NC2Y�4��r�{a�~�4�4u���C�4<����8��$���e	TY�߯�&'D�X�e�O��_��D����:8���1�lT����\Af"�mNk$��d-��<�D�('D���_�^��|l��c��'��DjN��Y"�? u�&���Z��R$YX|^4�[��j2X�u`�6�=Yr�m]�]Ǥd,��Z#>V�OxRݞ���D,�m5�/��-�x%��q]�=Y�$�z���lB������x'�@x���$�3�8�=4�Z� �ڼ�QY��qG���m��X҃cB&�����~,�).Cz����+ٗ�3��!`�ba4�-@�)"���9hz�W|R#��JE�drĢ�82�*�B�i/_�y:)���8fw���և�p��[[ �E�u:��K]�Q5hMZ���m�xL����:����$8��!z��$� �7���e����sp���h��+���{&u�����Ul
p?[D�%r[��4ZꌨS��ۅ":��%jW�P%�В�D�t�������:q��0?� �@J���կښ���t��4:%��OvyF7?�/�@S_}�̑�*>��]�y�j���̀�b�6����;�K,:�:�h(���<�jw����Nñ��eo}��MΌ�˓e�&�{��7��W\3xd�8��rB~p��?�,iO�j�ۏl�A�^�^s�f��f�m�C9*��4��O��_oO��Q~���&���y/���ѯ��p���%�Ez=r�iG��K��3���M��k=P1mz� Nj4|'���Ip���d�"���lK!d�rϳ.F��	ڬL��NXѬA�����[�Ʉ���b��T����`3$Єw]���<a��'BR#6�R;K	$���)��R;ok�oo��$�v�o�-T�8';(l�i�k╉x�yeL�����=_�f����n���v�ȝ��"ÿ�C'Gup�)�S�;|�LA�{��n�3d����-��=?"P`#��U6+��)pGʆ����Nc93x���ϟLݮ)�hV�t������p���R�</j���y�QOVL������ȔB��"�����r d�[�Vp�(Uw����������}�}]M�^�H�EqTw���qG!���.iĊwe�L�c�ʋ�{7}�2�t2���YyMc���ъo�:	�.��È[�]�d��}�l�EO�-���L��||�ؗ�~�+��x0��.Ԟ߃��0̝VzHE�қ0ѧ;������,��Ndq����jg~S�5n+P\�9FA�֖�?3��i�X�k+�iķ���ˁ�&�"O���|7
K�b�3�����M��MQ|B��̸+���'8��ěGO�����V+6_<fX ��s��"*3P�}LDRl��)K�V�.�e��%k0��yƝ�ȶ���s��n�z��3�}��Iք�bbs�8;�If�sW�@�(��V�ey�PCn^��r��ˬ �bU��7�7I��=�ݘ�=����������#1�K��2~�^
��KE�_4�K������~��p1���ެ���wj�㥩Yt�u�w�kKϝ ER�ӹ0����+'�6;�����j����j�����:�ttf���Y�~�j���P���q��wB���\?F���H_��Q����ɭ{4)L�����k~&N{��&t��:�=��WjY[�7@m����S~��.�	����ה��pE�L ���į��,���E���#}�R�p�L<��S��D�*�o�e@:�����6`�4�_'#����8<��O��b�Ώ͌3
i����p�NPV���i�/�e�gx?iy�4�Ø��C�`�A�TC0�d��{�4���4dF��&.G�V�z���Go6mB���Pu�&$�m��W�\�n�(;W����¶�&������|)O��~%E�{cp	�#t�5�zMǍ;W\����53��_[�B���&��dYD>mI�6�# ]׃�8� O2���هu��CX5ˈ��]'�����ԓD�X!��"��r�\�K5��	�o$D��&�̧)[�Z9��c����4���s�ߤN��(W�cx��;�{$��(�h�=�������T�=29K�W��9�r�j�Z�V�l����ܩ�\{�?�s�['�l��t�Bk(/�˿iL��6<~�U�}Գ��%.�؞��`��lg��?eRw� �o����V�M^���*��.��q��Ps���ь��X&xD��T �w�f�M& H�_z�=n�5^�}��У~�?�RB;��bI3�ˠ�c`�HT��|?�։("ǀ��?�0���6�J��7����3|K�05��h|ƴ�Pu����ODg<޳��P|7�[bi��5Z���1��I��t���_1%M���e:=�"2�����v,6�u��{��4����D�*���;،V�	��HMǉ�i_m��h���V�����̬_�9j�袙�YU�z�&� pn�k�|j\�F?7^3��*�;�vo�(a8���J��Y���wjp��qZ���Uk�#<��\i��b�c��.y��)�hs�47��kc=�����r�5}"������"/E�tk��+[� v���U)���4��ee� AM�1�w+$U�a�J��ei~�ˌ�x�4�W���"m�7G�!���c�k_@�ZK��G|�0��E�*��&�t�x��+	L᝷-ɀ�[�4~�.�z�í�H�.�l�%��i����S�[[ۃd���O3�uM�n���A�y�Njfs�;�V0�XS���g���G
�K+C��hy����a|����&�aq1=�t|޷c��4��#í�1³�`�3�u䢞9����ı"�we�9�g��z?*s�-���\?As.��