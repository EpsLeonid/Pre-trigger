XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��iswu^�"	��;�����B)���JCs��+�S��4�bG���u)�e�Fo:��vmWM��˧-e��e� ̞ز	E��K�E%@���6�_eޠ�ʫƠ��$���[G��2n��Q^��h���^��]��Q�Cl�LĜ=ˎ��K=@Z�"���� O^
��-M��ۍ�����<�nфH�3:o|2��\� ��ǹ*��7+�t�$��.︟>X��k%��2�M<�]Mi��]|�B���z~�Tih)t�Q�� ��
+�#ԡa��)�)בB�a����I�X���1aX��ư=�]�L���G�%���%����<��W��iM����H�+��}6�Z��(	д);���#Ɔ��@�U��p���+���u:�ٯ�䨜�Yz� ��?�ǎf�6���T��J�����0��
Ư"̈́�� �`+�p2�C'n���%x�1ܖ`r(W�dC����@�����6��H�&d��<Pj�a<���� y\\�L̳�b\6�>-�"]ܖr�|����!�&�!��q���Q^���DN��v��]�+�Â����\!Ch��'���J�p�\oP� X�"b�M!c����G�V��a86�n��>��6�n��1S�&�h�bm������t�g�������~s+�C���z�A��6�:�糆�{f�:��B��~F�b!C^�k��5m�&�fe��=I�J�p��Hv)�]o�?ur�!Y��t�|�q�R�:���#fJ�CiXlxVHYEB    5658    14e0�E	��9Zz)�_?�.h�q��S<��`x9�qvG˃}���D��Fk��gI��}Rڈrp��i�]�(���5VM԰o��w�Ҥ����t�r��z�l�d���Tb%���2����Ӯ8�#���P���~�]@�?�i������N���T��ALc��W�����E��z`�V���4��U�3���۶�Z�U��A�R�\t��� F���f�-)2�5!��QN{87F�8΋`�I��Z%��"�K#Q%��0AP�xj졢������"�b�M�����a���5%��Y1v���&������Yԭ�Tr3x~�w��P7�9r�s.\���_�����DT�x�w�ɢjř��X�nԫ����S�3��nG��%����@�D�XTTx������2�n�����BIV��&���~!{"�7���5���x΋HL���������!�R���Z�����fQϢ*�O݅�/D�����;�z*���*��^����L���!ݐ�~B{	FqJKl$���}���190g��A�����EΓx*SP���>D1.ߙW�4�g��4;]���g95h 6E�r=��w.��d)��.Tد�����/���˒V���&�ϛ��r��>`��i�>`�ǜ;�#���'I��^y���l�P�i��)'3�'Լ����9ңG"90� ���������.�����������D�+���C+Tɹ�[��[�&�����I�e������u���ii���Ͻ�q�^g�@l�Lu��i���6���]��՞Ӆ%�v�t�
�Ԙ�<Jl<��;�����.��a��_4��Q��AD��@a�d�:U��u�a�"����<S�����:g�:(IZ���X@�!�k��G�g�����c*A=�jH3�1˩/�#og�g���K��3���z���!����ò��"�﯈�Mj�B̿���j�ֹ4̗5 �RX��*�$!��䆲zW{!W����Q�K�+�ηc=G�(�J��y�Ws!����:Z���9��js3�Q�����
��_Z����I�U_g	�Ʒ��i���g&�	oxx�Ǟo&�mrJ���"��g2���WV�;�PfElj�����N9.�Lu���ҙ��r΂�̈́Lr��� 	��u[H ��~)�W#	Sh�U$Y*Cd�p��6xxk�ST��i�cSoܢ~np5qkZ{��,)�Mx!��Ç̛�9�J����=��yแĂ~���>��IBK� O�jVߗ��R�n�w���^���m�5����sN=����~���ƇP�X��"���}���I��W���務�h�]˦N�����{і��.��s�[An�W?�T�[�h`��*EΞ���g1v�H����^�[J.Rgrw�#[�Z7����s�-�^�<�iG��]e+!"^��NM�������|KL�e� � ��ܿ�h��r��V�0ޘ�_�l
a�0�������m�Wv��� _��K�px���!���o����	v��"6��VB��[J�ׇ&0\�w��؀G�l�a�	,s��LǼ�8���"��l�~_�nf`q�]_^;���Ĥ�zRd�q�{������b���&����K�]��� �aP�Zh�\v��V�	q]��O���N�K v��CdB·[�66D,-��"��PD!�D�.j��<�eI�f�WH��o�0�Q`�p�M��e��R���=`%/��Ъj¶��+�����+���J匟���@8�_� O��F̈́:���$�b6�h��x_3y+i>��t8�^�:b�����L����c�����P�v��<aii;4���u�x�)k�An3�:I����D��_7�'��ā�:�]��4�Va]~��ӿ��ɍ���}3	��.GuD|��-%GHj�槸��iƽm�-�2��n���hp���*ɀ���A\cY�7�y��;�enT��h��XC�|�Q�(\���>+'H(��홹-9`81r�7�
���o�`���m�2k���S��/+3)J��h(.�r@��o�����p��$g�״ZP�|�b�`O� ��!�mX�b[��ی�/�(uzz$����~+�i��f#�/�ij;9s�ȯhd��Z{$��L������Rv�CO�"P�l�uX���p.�gk���V�>����\�.����mVv����������h�S/6���ؒУ9��� �{j�SgK�Y'[D�Ǻ����c�cH���4�}c(��@�O����:u�-@�[�c��ڻw" 4�݊'Z2�&��4�'E���}�3�Rc�u+}����3y��&N��Ӎ!�*���>��N���i��7���"�q����0��"���XT��/ۼ@�!W��?V1,���
���5�_	�J|���9�V%�Z�W�eMq���w/����C�&�S ��(�zK����h��xǬ�wA��;�v���Ֆ����`��j�>����Ȧɺ
(.pqry��!�9�f�N�ρ�Xު�������p�)��k���n]�����ZR�^QV��?�!��Tp�ta�Gy����(��e��>�q�R�uta쯌R�H�7��e8��ȉnh5y�caP�M#�Z�,ͪ���8�Qj�{��ⴡ}[�ݜ��J~$⽐��蒊������x��¹�r���� [l���˷p'��[�u�M�0i�M5zP�Bp��/M�'���N���SU0�gq� �kqqv�i�u���A��Ot+&'xџ�S�(*zx�a����Q�'w�ճe�f�b�v{8��F�Ѧp��"�O����wAU��Z5�v��~�S�R*GP7��a���Dİ��du��oz��Ň��V́���î�N)3�vX��`���"T��㧅�a����
 >~����:e<oo�Ɓ����3��(�F���uZ���T󸥓�%iR��w�T���FsN�iA+<\/^ד���i2<P�����V���EW� ㉺��ƸC���M��1���%l[�+Z��Ev���n@�{�b�W�7��� 5e��iD��[�t��-)Ȋ�\�g��&��z8ݐ�jA��zǡ0,'M��N4>]�ٚ:=}��3�5� �D��k︎�$иULy���r5����o?�A�5{�G�d^� ~�G�c���u؀��Eʏ������Ǥ��w`���fB�9v'������w�%��UM�g�Kn���C�E;���0���/�ܭø	y��I��k	)����%��$҆X�@�r�![ӭ���)D�;�!�ES�V(Ѡ$΅[9�r]��L�a��I�����n��؞v	|fS]ؐ�	���f��M�}c#C ��U;p�0[ ����[���#E����	���gU� < 箟�W���):�\jb,�}��X�#a�GM?]�u�R�RU �6]�۷U�|dU%\�ʽaD��.j�*_&����bu�X�̝��5�>H&�H/�$7�2m������FVKr�P�R:N����e���|"���^�+V{�G�6�A�@���@8��E4���y�bG����X����X ���V��.Ѽ�����z-�\(���@+Z'v&����o��`�6:�U�r8�K3FH���,U�od��i����1"',1Q�
<�>T
,F.)��jԵ�Ε�	���}�Aj]�Sz�����Fr���Q>Ѡ��eE[����h#�� bYl	hM�Sz�ۈ�o�n}#��P�#<T�<�nf��x��۹�E4��Ԋ'm'Qj��Ʃ5�dGu��N, Y�5}gGv5��},��Ug"a�����,60k�RR:�)��-�j�i�K|P�-�z����ɦ��Rskyk/�	"�!��A�_�Ժ����=R�E�@D�*��sV ��8�f�H9�Mb������^H�lC���������?Z�zu��������	��ku}d��U���\}^�?�B����K��U!��D�L�ݔ)ی��nĻ�yd��Kyw�	&��d�5�i"P�"@	Uv1!R�����*�$7ȥgc��V�uH��z"Y���9���=�~Uq���`�(]�{��	�����Ų�2���<�bKu�Ѐ9*	!�bOT�7���X������ZS�kP�0k��H@��߼�cYF�R��fV`�^HLȤ)X�$�I쭑���(!ӗ�ꝟ�S��򴱄X�l_�<���f�+;UriOo&����:B�"��V�v1w2�i��27���t���k�T�
!�{p��T�E(ZR���x�D�G�[��M�9%%�X^#J��mb��S&��T�n���*�hxYȀ.���Ph,�5/o� �vYse��	Q�Zu&;�Vw;��]F8j�Ej�g�R��PF�ޔ;;d�<IsT@F,<�Zf�B��k�\��6؜���,���4�W�G�|�c8�\���l�:͹\M�⫁���n�<�W�SHNޞ��Tf�4W*gf���l��=}E��n���wdfM$�"B��n��]�̝',>0� ۰�@��4����^�҂����F����`����󠚛���� �����}ޕ��� ��-�z�hMd�㝭F1+���ɼa�z���,��]2鿕�8�[������(��!�7z�I��J���r�.����(n�=ܝB���\�$ �g��&I�gy�}�oF��F�p(衒�EЖ��|}xu�y�6��������J�8�>~�|�Vi�ks�(�&jpضҰ���x����<�n�`�D�E��	���D- ����+%��Ej�ʾ��I�k�L�z���<+VD�s�$���4����D�ND'���E2��ƂX�ތ�p��}���\rF/=�>lV�$��|��mBwe�D������f��Y�����K@o ���=�_�W)��(�����_�U��	���_T���IW�a,]O]�RO0�,����`�i?��7���ŉc���&z;�@}��V���-p^���l�*0��+� �h"�[.��Z���;�A�u� [)m�5���wU��~A��ZG��dD0]�g}6���6y���_�4�L-�����=�ۨ����5����TZ��ϧ�;7J8y�7Ɂn�<����Y��H�))i'�l��g�xz3�9��m>u�Ha%�Uho�9������Z���
�m\�x�g1�p��u�䮎�H\Z~2��H:Ŗh�:�:Z�}.��/h����/��və-��s