XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ߎ��fY�75�����Xʛҏ	��߷�~�s�v.�>���9��ȯ-�N�� lY<���(��30U���'�_�U-�K��GAf���#���ٙH}�/:�F��:~c��7�ViZ������<Z��N44.�#WOQ�A����%�pd�y	�A����~&Ì�zUƜ�8GLw���'�y���Pe�h6�"ܳ6 �J��h{�~yJ�ّ�K��	G�F��&+�^�d�G�$�a��&T�A�a���z��3�.]�-����c:?�+��Z��l������jC�PE߃�Cx���ՒZ�v�pk�6�;5�I�g)�K��d5pڰ�iV��D�I-��SY��E��;���a� �C�uZ�𖴣[�����x� ҩ�֞dV�Fb��[ء��!0���f�����wJ����8E��Ѧ5��B�kC�=�Jf�[p��tQgYG���qA�)���ɬi��:ˈ&�����{�r�*��$�]S�{A�-D��}��t�u�A����%tU�n �Z��\��z���&h�)]�E",�C�7�_�T�����<y�y�Я�0�xO�K:��С'[����rޫV����0&��d(���&��{��L�|������+t[;���Mu(c�%eL���e��D�Z?A�|n!1 2��au�Gr���4�P�gFf��p(���:���F"�<HLM��������}g���-yY�5�~���]���R�$>��˴#�8Y�#XlxVHYEB    1e12     920g��11e�݈
X2��.Y�R�Ta���ʷ�y:0O
H���OK��r���.�aRv����rz��U��m7k�RR��6i+zW��Z{��U=M���>�ʩ8�Y�Q�\�B�^C��r��(,���izAg�7���G�.���W����  ^���Dt��E�CSï>Hѹ�o�59�"�h}�#��Y����%����~���5�ϴ��4UD��^^;h0��4}�&H��&bkC�yU=�������!%N�Hb/*�X��	9�������E�?�VUh�*�Ű��ᙐ=��x~�7S_��� �8�	�#�e�*�7d�KM�h����Z֠DR�*���������=���(�Ev���Kj��]}�_ �2���z�*QϹ�R4�t�:�,��U�a�^.�?���M7��N�M֎:����ü�i@8t�gaJ�u'���p��Ziл�,Q��˶�籬�0*�pD�Qq����t1L}��D#傖v���ڂ���{���Ɇyj�:���(�FBM��O �;�8��:p�厼_��"��0����]���� pw$s���e�N-����<H C��#��q�#�=z­1	7hf��0$C�o腺K�H\�[�Q��6I��3�S������U��L�x�U5-S���[ڞ�y�M���Bp��&^-p��N��}�#e����������Y�2�k]S�q,Ά�h���G7w~Kux���
����O1�W҉s�b@�ar�I灍L�3���FX?w}��5�b�Gg�d'�>'�5�U��FX��2��8x�/�6���+�4��>7�6�����z�֗  �h��Ӥd.�&�Rm�3���|�w'���.�9u�L��0�{[�mgތ���C�[�}�U�����[ŧ�i�%v�0����AJ8~�S�i��3�⪤���懸��Թ�J�^L���u	p��D���wۣL�Y\J��0G��&?��p���3���r�8�Î�)(�]��[����/��t�`�Ý�bEf� H����IFؖZP��΁�4�|�,f��Ȝ��Ư��/=�J�S�����l�C�:�.��=M~m7�m*�d��V����}����)C��}�Nk�2���_�����}A�����kk\������
��g%`d@��V�ܒ�x��ԚI&�ʡ޷6C{q*��xV}9<����IY��ŏ�R��n,Q�Oؿ�R'������?=��߲�;iخ�&my"��g'-����S��ӕ�y�r_�((��:���7pV�-pZ[g J�?/����P��S���I���A�{Rj��'���;)��Cf�q��W�!9J]�'�WT�y�'���HM"�>����[�����n;�,1���!�\�y/�Vf��
��Dh��qF�	�	��GT�x��A)e��J�U�//��F��~���v0�$O�ǆ!�N<����Y���>(NLJ�f��	ɽ���������UE7 N����S������$���kf��Q��pH[��1�Ĵ''�>����u{ޓ�'�JP�@]�H���~��pZ��bNO��;��N�؏S=�%@�\��4������ ��J�^���jc�������ջl7rӬ������ׄE��4Gކ���#p��������{�*q91��92J�Q5]&q��۹�@@d�i�nfs����K�2o\�N��� �`-���h��jd7�̛�(P���!����`��MwQ��y�l�GpO	��g,l�S=�����`�R���bMg"Hr-�f,�<M��[�d����6�y�U�NAo|���%�`�}��C�%R �:?����7u���������lJw9���(�p��@q4�ٟ�b�V��uy?!��o�,�O�"�@[Z�?�50��&�L��"g�d��,�k��cby�hE�d2�7�Z��V�	F>d���Ǒ�������f�j"����DV����,��':[�K2�:nZ���Y&6Ž$��E�a����k)��O���a[�M�G6�WQA�8��F�v����B$�(��!�����Q$���e�6�8�??��C α��p`�x�ip�o1�n�o����FշjqM��\TWz������S�����K�2L���52��!�����x�'�`���C�3!�E��:s�B*��P��`ܿd_�ӓ���%�;��i��TZ��8{
�W���c�� -f!���P��%��$�5��G�I��,� �qFg�wm�y�\�������E%9�R��sd:����I��g�rT�r/�BCOKae�K