XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���
Q�I�ޟ6�	=Yς�)�`d��*�2E��D�Y-�<�#<���j*�A@'�_m+�y�(,1���
)( uq
/�^�}�r_�����u�V��_o4����C>���y�6�4#%\�����&��F��V�C1i/8�8/�dc⧋��<�.�"���¡9h��)A��રՍ
�,�s����U���[�q�QL\ў��ȉ}��ӻ��X5�)[W���i7�x�d쿂 �<��i*�X�>I��K��y�_K
p�f��y�gD��|�5xzy�K��	�[���C�\���'^��x�7�j_�k~B�y]m��'}��Y�${uB1���N+?0=��ޯhԃ��Cv��@��jc�O��6�!���r����oG�ϑ���LU��<�V��%��p��=�	�ϙ�橒��e8��z��|_3�2�,I�[1Q�BK���R�qG� �CZ�lD�E���)��3:~-�#�-M���-�ߍ��KS�خ�5�Am��ª��w�)\����ץI�eL�;�}��Ȇ( 'L�N>9L�Ȳm�>�;���$\��7:�4Љo���z\`�;�vX9$Ը���پ�¦��م�vRnY�i�W<x'�y�L_�=ת_��iĄ ["wkGTk[�2wI˭��4S�J=���J�ț�ʫ�>�|eC�5�]v���pQ�=-�JK�DY�H�K^�
q��f�C���9S���N˕fcQ�ۈ�~ǵ��
)���c�]�{�h�Ug��@�#�T�XlxVHYEB    d81f    26f0�j�Z��H�}�Uw���ޏ�\���y�<S�!Gn����7'.�И�ya��כ��a��夦�`LSeR�������|�%�����$ut�O#���ߌ1��f]�9f!<-|�y��5?�lk9Ж�	�Q���*'BC�-�uRJ_(�(Wp�p�$�� .Ϛ�v�+=��p��Lբ >C��{��W�&�P �O��J<�?R:��a8�!� �ri�A��z��o�V���ó��o���"a��X��,U�:��hV@�)PP$�܁��ga�%�3�H{��e�YQO����9_y���S����T����=I����ǭ�;i�2��z�:�f��x<�[.�@�T��W'k�Jie��υ��t��t�3�K,8ˊ�+e�����Tz��P�_|���R�Uބ��#��e�B��n���s� ��qT��0	j�ak%q��1��X���͙5���H�cm�Q�*���Аd����S�I�8ZqI#b�*�4�Ͳ\���$<Y=O��)=��W�,سrS1zx�R���1��)*��ۤ9�y��Fw�$��'�qh�#6c�[y��̮�3���uu��^C���D�)Wm*�k�n|U�$�����?&�4���%���%��?�+�:�'��³�W(İ�u�]j>'���'��Rc��Q�i&��w��yOU���� 2\�3<�T�c��"C"�˦�6��V|w��6gMS��U3�y�����R�r���g�/�����&�n�"���Y��&f`��=�L<Jl�P��id�%�����eP�������0�/is ���P�DKE�2#��q�ˁ�a�H��b��v���[����/U��Br`�k�i�S�yT�����O�q�!!{��G�Jg:����O1-"�S3����լ�;����w�pm�w߿?BiԞ\�0�Jqo����>��[]}c�N�w��s�w��F�՚WrLU(ҍ)��Y��m�X��իݷj['ѳJĮQ���e��;-[=�)2]�ETewЫ�[��R�u(: ��/�q~�5�Z �ċ�$�E�B:FQ�́~����^]:iK�X��Yq��)G���G[�֤��9�%��v��^v����v�������#;-Q����⽀���l��Fl��te�w����G^�Aq�sQ���5ݏgy��4���w ��4����_��I�}���"��#[���m�����4�X�|��ћe~�^3Sy�S�ޑk�S�ϴyȨ8���?/���ԖHn3�x�2]�����<�'��������R�ד��~���Wv+���X2B����j8
�76����n�T��3f�=�<GO��pa��A*`{�o�>!*��#X��ұ�>]��4#q���4^'�8�7�?9�@p�].r۩�BE�?:'O٢k�����'/'��٫bA�q-n���>���rjӦh��T�iL�G��&�!>x�~�� :d��ZM�jF��v5�W����{��Z��Qﳕf� �;kf��)4����3�C� �Ld�� �4���3�.L�K�����@܆��=��_Q*<.r�]f��)�+�Q���`�!9�Q7�>��<jM�X:]��t�t��>q;��~��;��c���g0�������1�����5� �\]#�0�;��-U;$�������{�*����Su��پ�h���w�<����8�~�w�9���[�v3���{ �3� �S���sĳ�]3[i�C��,E`���W浅#�fZ�x��X���Q���hd5��_�W`&�/��5�A[�nDP�Lo�,����*�˙l%�Ӎs'~�����$f�=�Y� C[�X43�Ӝ���^�J�$��x�m)�U�oӔ�g�����71��7�
=
u���RǕ��x�38���>�'(#O�e�ɣH�L�j�x]�ߕ�A�^e�ؙ�yGs�_o�ܤ+�O��� �}��.�2U%��d/��Z��H$�jp�,�VR~o�ݝ�R9'pR����i��Ԍ��}ʭ�P�H�
�:�|篂S��|�swJ�֋
U&N�w�Uo��?J���}���0y���Oc�gn0y���Xֹ��pu��<��t�A��e�Q��UB�G���r��_�#�����Y����*6�􎙦�f��̙��\�d,��s��.��9&з՜*��m��z��U�!�����!���៣���o���࿂�Q=�4����N2$Ny�YJz���/�����=������q(?ua��KG�r�08^��"�|�r��IG��s�Y�B��s��MfQ�۠!��2��<E.�A����ֽօ֥�J��ryL3����5�h�v,v�t�gx_���w�0,�χ����$!�iiF��/U��m� �
���BU��>���E��_�p�`b�q�:l����EEy�k~3-]c�X�b��[\��.��'L�J96��xd8i�y�@K,�U���	�=�4��h���1m���7Q�8|�,y\Q�s�NTd�ةRd�<�֓���{p�վA0T:��*�%��e<���Öm/%�Z.�7Oa+�����EH���� �A?�r��)�YX�(�в~4�?�e�E��k�*c3(~���4�P���N�-NR �%E���F�;S�Nw�+6F�Q8�>l�t93ٽm%�S�2���d��̡�k�؜�»�{��Wz.U����`��NU/@6NIG��)��K<Q�տ��KT��+�,�y����z;qt�K���o�����t�c���fS����kf���6���sG$7�B����u.-\8�d�T�	����DYfA�j�T'83l�[wUQ�d��я��y�2��vt��A�<�e�4.�7����)X�/b�I�}_��S�ZЅQ�9����%CnظP=�[�7��s'v8Ffea6}�M��
s8�T!��+�^b$�%0b��+�"(����X�`.ayZ�튂�8�;�x���D�pM�oAw�>q���R��o4B+����G�fռ�q����UMY��Wp*L2/j����獪P!����I��SMң@D@���b?��kΐ4�Z�W�h�Q"k��i�%��$t��JC�V��A��=�Y��H�Ι�>I�k�����]P��C�d6����b�Ȗ����]��0B\C�i��'���
?��	�s�z9~������D��^U��y�"��po�L�	p�m�T�RW��&��M��t���͒yV_?[�}q�G��[��ا��kcZ��GΣ���)M���h+cm��MP���BY�C!x�rd�r��e�qՇ��M"ݼd�J%	�uT�����J���>����ь�z�u��s�in@
�;@�c0w7sZ2<4$���Ë��Pàu�_�q_:5k=���8W닪L��l����������I���0��i�!�nJ�+�"�|r�9��0i�v����� ��6�5r��S�؄����t8�r��܅k�6�1?L�V�Ϝj�9!o�3�8i��b�+�Տ��� 2��49��!�A��E5�=һ3K����V �I���CȀ��7��e��`b��G��&m��6�j�0�
����8;��d7~.��c��_�&�\�P��o9����n��8����&e~Y�AVI\Qt-	�Шǖ�3_(,��X~��SG{���vB�[*ή�#ۃD=?8��tv[���x�[�=!�T���� ��c����P����ޢ�����I��:
<T��_d��1�ȦG����2鳛���$�-S�gG��#1�ˢ�� ��R��!�$��s�f��Ƃ7���O-�#�%ON -Q|b+E��̇��f��5�S�������:8&l�q�ۛm��&YT��?C�[�!��$eK�p� cb �j��ə�������s#���v=��о*���x�󵷆Ǣ� �I����	@�J���U��W��C�fN�3�� �wV�K��y�������n�g��͟���c �χ9�@k��|��}V�ǥ
��9
�v�����yEbf�نXֺl�t(<�r�r����0���鷭��g�p�y��� �9��Uubee��E���8�0~��Q��I��GD����p�=8��
X��ꟗ��V����
����P�JYU�z6��|e?b��X
1���Zc�.aj�i��J��ߜ ��}e�Ô�ŷT/J�-��J�ي+���&�n@��A��H)����?w(O��F-��RHYm��u�,_9��8�����R6z_6y��Q�jF�^\�4W
���0'��3qn�u�i��oS<f��������ޮ`��>��i��T �!]]�uh�t�Bf/ɾ��9	��߉U��,�U_�h5��}Ǘ	=x���N:�'�E���L�Cg�[b"YN�*��¨Юt�rF��n�Qi��4�u}���rY�S~�<y��"(:������@~.�`�bD"o�y ���Va$�5ǗO�W'�����G\e%��!#���xso,x�+����6�H/u��We��o$�Fr]�lɌoc��g�I?d���НH�</��s3� �O3uP�V�r�e���	�#�ʻ��k��5���})U���'�M/Ȫ����N�n�|���/V8���
FG�?�Ӻ61Yw@ ��<Ó�k�A4���俵a8�+�ES1$u��VP)�1�5&���P���y��߻�@�ٯA���M�#/B�k���a(h)uӹ׾^��)l�4�I���f�Gn���e@D��]�0���lwEգ��r�N.��R�&�g�{��iB�̥/$��S�)v�0(���,T�U�	`I��i��6D���쳸�b�L�<���ψg�.�*������r0/�d�Y�S�^B�+.�zc>��2��,�®7F��m5�)]L���i����v��4�Z*���Xc8�G��Ά��W���Nɏu		$M��.)s�+�G�M���	U&=�=��F�1%��P�|�t���L���՚Yª��q���)��!?�2�ǂ�o�q��b������r#��xB�u�M�6���[���z#ӈL��͘ޟ ���[��2�Q�{d�c.*ѰC0��<B���6��,�V������QO�;AJ7)�M�w�W|�ƀ�!n�/�af���֝�;�a�q�.�r�&�uy^KF�G]Y��`4����-�x7����×}N���G�v&J�0����G3.����/W�yo%�,����.��S��rS��_���w� �|;L�����ɏ��Zġ��8��w��7)P����6��p���B��׶8�X��ᕌ��Q�)=Eo_1���`4vw�oLr�%�yy]l�4n�O�la����h3��h�[��:_��sT��"����Y�)���bL1 ꍈ"�0�q�5E���.e���p��r��CfggÈ���Lb�����Z�GO5v(��U���@�h�	x�Y2��3�?��̒�"UDR��ѭ$�[D��w{J`qҀ�R9����{B�%q�x�9���<n�|?�\ڥ��z��',}E2@� ���o:����m�a�]\�dOS��^��e�T���7�'�tr�!_�����P?j�ldڑ/�O�eG��J_"�n\����z0�p�~��m�j�[y��,�����8��5@"I��n)�S���!�c��͘���H[��-��2Pt�o��&�v��J�q�ȱ�����2�cߕ��2(}����"�-ޒ���4sB�揗(����ˣo �?�������_j.f�׋h�������0���W����<}�n3�X�cF�G+$oʘc8j ٶ�^���ç�3�4�����=(�±Ȝqk�#Z�X[��	 m�1L$������J�qˤy�#���uQ'9p�:��`��bSN�t��2���cPKJ֑4e�X���3{�qs�2I�)��������S�(^�e)_�T�PTV�}�`:Zg��H[����9�����h�.��ݮ�<-�a��n�ƽT���(l��� �6䦾}vkuC�4�� ����u�dz#}����%�_8Zh����@I���n���o[�g����SԴ|�T���-U�������Ҋb� ~G�	��]�tp3p���'g9:���r�8l+e������'��ɮ���]��*�A��I�%d��#  ��lK�^{�T\n�9�E[��j�=�d\�?c�H�7����`���s*�P��G�<�1/v�Njx]�u�I��d�h�T�)K:^������WsG�2������b��A��^ϡ�nt.��()�/wb 
9�}�u��>Q�.g��^�>,�������v�&@�y[@&&S^�e/eݝPp M��P>�tׄ�,є=܄�o��� �N�+�jz�Üb����E���}}������g0�7�0.�O��V3�4@�G�����,�s����nB%A��|�}T�>6ǳ�#��mZ�N��[�[<	��;;%.;�i�Lò�ɣ2�6_(��o_����s\�?��ʠM֠�t��;ȢL�KB���z�����<`��m��ج�ROA,����&Z�ֈ^ʜ/5&7R��4q�'��ŔT��r�Z�ڔ�� ҡ_��f�aY�f�'�Bb�h�ն4��ERYyy���By���$�@}
�7aӔ�w I�b�?र�P�L�8D��
�������vA�/cbB����ꕴ��]�Ƹ�9S���'l[����(
�p����;���/%9�q�Sפ) �h�m��
�D��}�+_��K
�K1��_ܪ��"��bIw@K0����������R���Ĭ;.�R�@����j�(E�׹
��xÙ�����IV�B�ro.�} ��<*=�8gK1�!� .��"�v5ߣ�N ������74c���
���cW���4ac�+s2�5FXAaa<odAv�-�s>d�H�b����������͢Џ�d��E����CܜH��co�	��\�SUC�~����f�R�f����΋�ӱ����̬d@ր�5����#�4������pL��R�ȃkJ�z�@	O�	���`I/�[�S~M�l@&S�
/c���{�0)<�8)s�_	��ᒔM���1@�Rό�<쒉��^JF̹S�>�j`� ��.��9-��ptq�K�F����m���Sk.��g�xāb7r�����Z;O�;�޿	���o��{w��|Z'��bp1syi�ꙫ{�_�+��5��ә�@7ZcO�HGꂅ��CJF}@b?�gn��˳Bp�Z���p��b�� LbT�u�)i܂��m`RR@�f�w�*�΃���}<�}e��&�L�|�nyR��z^�TL�R`j�2KbH��q��Y�z���ǥ���&S)�r�������K���6�3�1b9�̅F%۷���0
���\l�l�a���x!���Lu?6�#~��ٛ��T��>r��Ѓ|b�¯к��qaM����x2��Z�Ղ}h�Ù���˞>����i�G�#�;�z�t��=x���������=uUZ�R2*9"�$����ZJ4(�Y�XSMT���W&�D^�l��UʳSg\�$�?�NZ�҅6I�/��BI�%
�_An.���ΠC���<�۴�9 ��hW.�j�%�[��23>�S�wϷ������j�$��X�����/�����#�D3���	�d6c8��/������џ��4/�)zy�^�"ٸ�rW�7/�M��ɜ��A�iyr/�� ���u�^�\KSQ���%˛����gR�jC�_P�q��'�jӷ?�^jVSk�L#�3HT��B�1Y���Z	m� ����1��A�����$~[A���=F��E�u4���of� �9�ıO ��݁_�<]ҏ�WG;�E{xs%rhT����OqE�J��[,�oa�QA�iw�^I�Z�&��)�,"x���Ԫ�&/w���V�j�d�>�X��>P�^��t�i���O~X���"���_.*`+t�:�"ɰN!��jх��%�@5v˧��5̙��Z�n���4��&Z��u^����#9W�
��+H7�}�^��t��I�C�r��c�6g=����*�J��=��盃\#�c_��vbp���H�I�]�@��3�r%�%;GԄ��(���on��L�\�2膯�?ѳ�^�n�͊/�����Aiw`U��Ƨ=�*��X\j����Q�(_É͸ȅe��1��Mp�G���p���]TL�Ȝs��"��]9����S��%�q�Li�+�dp�A�0�GؔX����7��vEJ�I6)F�wa:�:��A�{�B�,�Ĳ�1��%<CZw٫��̑�ݚ*�Ɲ��ʁI�G�J�2��Sy�A��74�����C>��a9n���;wM~��D�Z)1��f�T�0t0y�V����]����!�b8M";���G���a�rcU���Q}��k�n;���QQzQ���-ڭ�fE�UN#- %��槵�9NR�ޓ�)�"�s��,>�L$Y�_ّ
�Q%m*9�D87��e0>:U�)�1�t���������Vu�^̭-YC�~	�q��y�ڣҺ��:�]\3��5%���Q�^�$)b1���G��M
�v�'6�]��A21,��U��GW��in)v��-����i�LDݰf��t�)M���BPf�,�1��!N��X���*����QJ�A�	H�PP]D����v��"�zW��)Gn��ێ���3�ӵ��T�/B��z��W��c0 �O�U�/�
��ץ���*Ŝ�mz�{�f���ۗ����5`��m���h�s��ZǞL0����*^��9����Ѧ��L�/��T�� �.�l(�|p�z�K�r� �P��3tdoBT�Tr�c��Ȯp�p����N�4�'�^/H�P�u���o�n��^�:z���R��[��|A�����2�W���Zt�8�o�KV�յ�\��k����UHѽE�#��a���@k�F�|��۩rSt4���T�cΣ��:�a1|�X�������ϳ"�D���
�lX���@���,Z&�K3����\��C�����!v�.��H�'���)��Ӣ�'e[�\|�9'^�ig؛�dg�".&Lk���"f	��Hi��6-���(P˨P���I�L
=�	SIL?��#� �j����]P�K�:�if��~��b˥�o`��g�'Ri�h�g��A~�G���d0z�a@�4�2�4p���ϣ���,�-O����E������o�h`��U�����A��/� YZYU����H�4T�$B·'��XZ2<]�1�2�+�ҩ@9�����`�\�w~�:�4l���sB٫G�3�@�Z�Z8�D�"���+��	p���O�W����,�R�*����м��{]����a�d/-���_�?�Y��������� 8���1�޿Yn�/�x>���vy�Jp��Q�ڟ�����=T���M4����(�ت"���|[/l���?���QUO'�ҳ���$�4���� ��n���y�;�F�x"�CS�1�))A��O�5�F�[m(��[z�^x�?[�QI"�Y
�.�E�$�R�iYRh�oc͖5t������G�F6��`��D��|�Z��9��#j�QG���s���Cei���������9�}����U�'��� խ��P���i #��p����,�:?���L����