XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���@���&���H����
�3����Q�,�4��$�X���9�U������a<���Y�[y�U2� |��\	Q�yW���������_�i+M;u�j��
�QL0�iP�j��Mv�Q;�ke��8g�D�%��X�� �� �V�v�x$X���_�c~�����,�H-g���O�&fn��Ɖ@a���e�.c{�S'�����u-��m��yy��7om��w�F,�D� D��o�"�:�c9��K�'�h����:�Q&9���] ���ޫ���8;���B�8�w}�K�-�����Z�[���A=,��ײ�/��v��X��dbP!��w��x0��$�5����] ��t�M�χ�!���T���0�;�'��_b,�nf/�w�����0eF�PH�4��RM��]U�+&��R6�)�G%�E�ka|!��˜A�ߝ-��X(�D_����D�!�iV������߯>�Qҙ�NB���޼U�Ș9ZUBA1�WAd�y»�z�]�Y$3VpD(4	��"���ȃ4��(s��.i��!(Y����꿞�>s�����p��G�歹LY�j�����Q7�j9,d��=/29ʟ��
7&�WvH�}܍�+,���Z����4�'��!fM�%ǚq2���fȽnk@���Eb��t���xk�{�?�.�~�L�AF�8D��1��Y��T���0-ڑ �oh@>��F"o?�j��.%�D{���t�+G~kJ�e����XlxVHYEB    1d59     8c0�syK�]��f�]*BZͱ�*�f���FN�(��N���+7�]+`�]L̳��F ��]$�<]��>K�͜$�ZY���*��0��e�+�'[6���C�Y���d������� V������}?\��Q�6��6qq��L�*W�b	��ݙ���jM�}�ս���r0`�cv�4��Qʾ�vN!��!ք<�hi�?�J�K�a�V�O��t�0^(���t+U�yGubr��_�<h��g��\�B2��+Z4#������LE�/%h�^� .- L�:��t��7R��2[�B�$��_:�9��E?�����ōI�[��>��ش9̞���'��xE�L�b[�������H����`�����C�%?u��n��+ȉ��r��+����+'P��3������B)��qZ�8�_�\^8;��	�h!�*�m��;��[�M;,�`؈��y�{5����j�,��1ފ+���=���)�8�A� �u �:�&��H���� �W�͙�ꯊ\��a�L���ȉ��ZjP�/t�_d�]N��e�w�lS��ذ��zS6�h�릌�l��^���C�;�u5J4�D�I �E]��+�C$|�5������1��c	�dI�p��&Yk�PN�d��Ig���+n��4g� �@ԉ�`��!t�t���UJ�h~�H~"�M"ݳ7[�E�L��u}�<���mvJH���\�D�/�T����|��g�.k�@ ��ȭ� d^�T�e��A���̢�N��pJ: �������%չ$^�ywÿHJ�JF,䝡��Auy�t�7�%� <*��H:��ő�1Mق>Eq�����qH�¸��� #�iSn{���ր�3��$/n���:�d�{*EQ���	+���C[�~g��訁�s�)3'G�#���{g*x�NV6*.���){( ..�.�, P�&v5#n��Ѝ�Gg^��%j�sb�˅H�]�s���л"��՚9<h]Z� &����Wk�_��Eg��hy;���/���q����S�`#�e����o��֙�T����������\����w�D7� A�c7���T��*���ػk�Bk����Ѳ�9��Romz�Sy�nd���r�^ ϱxm%�&��� iHj��7_��e@�M+��<*}\�l�q���
������X��η,_iM%L`�����s$�ېN ����(8R���ٝ���r��8���6r^}���5�ih��KΗ�x!�1���@��W(�L�3"�I�e_5�t�Gq�����sħ��70�cg�ڥ������@4Ɏ���G�&��<fhb*�����PJ��AY�X�����+3rk9��w�>'��&R�*+Y&¹�|A����o�*��۷=�-(�%9�\a@(��q�F�c���/nK����&UW�r$��l�>a�Q8`ٞ�v0q�t`l���|*�;mgB{���k�k��I�ۈo��`#��Ϥ��Q�vo�G�P�����م�������UNv����x��Rp��D�y: �׮����	�iWa�c�(X�{��TK�hӨ�t�f�]�D�B�#J�]U������^1>I��nU�%n5qu��1#���r��h��_H&BP`���ꉼ �����J)�5���)�9�*�z̄?Y�L�T�btӕ�3E(3�lט��>��Xt^��F'�8#��5�1�τ��۵ˀ�n�����-yK�(�2�<�\�%�$�[Rv<R�ߑ�_
�J�u��W�ES:p�y�@��wv
������	3]I��\�-wy#g�X�X�H㞹�
\���t�����
M�
�Ip���c9gA�)�\z�~�A׭�}=1t�0��8|�J�>1Î� ��C�k�F�T�V*(��0��������JI	?E��9�3T����?�뗸��=�#H�E���P!�t]���Ɏ���t�I�/��[���\�J��Ȯ݆�%�ؠč9!��[���h]}��0���E��k�9b�Sv�{@���R3&5�
}1�X�e��,�g�?�u��"����������Ӊ�M5���Վ��R��x�� ց"D��\�.م�*�����Ô��P?]@{eA��������q������7t9� 0A���\�c�1R�J��χz�Kz@%uBI�3#ӯe��0��4"�ݩn�u�B&ǀ⎪��