XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����[-��,����G9MK�Qy�"����ly��ü,�	��M2��؛B%>��6��w%K��\U���3�ۢ�S�[:EJ&c�ةDc�5��꾡ͽ>���E�ʲ$= ��Y~�6�n��� �Y}�p�S1�A���<Cv{ ��_��f��Ͽ�:���b�B���A�P<l˓ͻY��,!��&
ڋ�E���w��V\g��Z���ΓJ^��>!�C����Z-��n_���i!�O�u�X,�h��t`;���K|֊H�뢞�*4-���c��!�#Q�?�8ן*��;��i�rK>��/3�y�A�(���#�����
�&*q�Y�e|j�nt���b�ҝj����4�`!M:�!OnTƞ:����d6�5�B��A�)��ã�vb%o�Q��q�������=�/���]�F �Ρ���+�9��k|��9G�ǜEjHV!��6�y��@|�]1g��rZϣ�y���������2�����p)��wG.^=�����jq���ʭ��>?d���:Cgl���bh9
{Y�d!�"�qh�H&�w����J��pv�S��",�Rݝ�s��Y��j�[,F�5�ʛ��(x�$؞mjt@\!���<a�4�x�<�㬏�W"�L�m�6";�Ȩg���%F6|�]�
Z��)Q�7���6�g:/q�CɒT��-'��U<�j� ¡�ǯ mLU�	���'C����R�x� ��.p�{.]�e�Ƽ�/RQy�O���>p8De�v�73�p�v�h{��BzXlxVHYEB    4c95    1190B̟��\�]���"��sw��mΫu_e�����~���1��,���:a(����f�I�G��
E@sg�
gT��-�t�Y$�A���|���Q�ߖ����5�2����r����BQ�oc��?E���q��HXX����JrtBv׮~���*,��V/'S�� ���ED�7U3�z2���N�x�v&J�;ӕ�,>��/ϒ���%�^/0r^�}tN���Ӣ�0%!1p1�311�|6Ն���Ko�v��5˗�l*8s�0rG�����.�|b�Re���г3\h�������E�?�X"�������Uǿ�=�;��rC��Cr����d�#t������J}g��0)�r�ϲaYBs��̔-`��:m�Ky�]nَ�w���SXݜ!����р�܉P?�Uk�%a��p���6�WM�I۠4c��15}���Z��襥�ėkW��Â��"�������B�I������x���q��~�{��o�Cb��cA�2L�[��7a2�;6�6�/5�D@�aZ�EE�0/���?g��)�mJ�B����6�Ge"n��6����~kBw�Ns����_bF=V�vU@L��b)���g���+�"�ё�����O��*e)	�hc�23*��w�PahW��ک��T��ح�b���/����($��(��i� �n''��%�0��.�����U�����DfԉI*,�T��{֒�>
��*�����l"��K`W�����\�To������`�uW�!�P7c�c|�t-,;���#?Aphɱ�$��z�$��)����W�U"��@̊}o=1/o:���ex� ���9a?�����B���?�KH[�f,�����F[W���K�&�!W����bw Jӓ[��t��0M��&=�x؃N�Q���jѧp�xؼ�c7�yR���hQ��Y��,vq�To�'=��u+�'�i�H����=���@�v�����%)D�����A1�cA)�6���@7�P�K=8$��fYP�ur�9����&ڳc��)�7e{C���l7^����C,`��A��h�,�#ou=k���i����F>�_��ܡ�9�W��Y�7z�s,H���{8��Qw�.$#��\�g�Qv�n�Iyj ��)��y��q�CxP.�t�"e��{�I�S����#|a�ޒΞ����W:�l�R6�L҃2�D�al�/�3�(�>�yd��\2�P��m{�h�k|'���Ԯ��w��t�D���yÉ�J�`�R���A�}@�gչ|m�<���S�,���~|g�	x���G�ëg�ͅ�B��,_�ա ��T����=vǺ��V$�ƹ[J^VN�\S1-�V��u��<��sg�(����@�E�lvbB�?X��F4��/�\pӔ]�? ��-�eV�+V�3�"� ��h]�h�	0��a�K&r\N�#ڹ�B�(0�vklq�3�-�RV�ꄛ-�#��h�c����� �⽘�z�%���@�Y��t&^�홨i�D��iU�N�VƬ�g0��lH�����	�b�����-A�>�ϳ���;�Eh�b�X���M?t0K���7Vw迼hZh@���m}�ds��#3�pl���P�f�����`x�?�H%�-~�j�5/�/�cB�V��s��3�	�4��g�X�ZN){ �#r�k�BxQ_���G����e~�8����hZ�𞿀�����B.�o�.b���H���a��.��X�l��ói�K���-7ЗI�vf�;:Ĺ<�,'rA5v���W�8Z�C�~��jll���p]~GYȬ����A�/��H���\@��@~�z�w��v�O6(w��Q�!�!�z|ڍ�m;ث)������e���\Г]H����C�E��u�9�]�����~Qĸ����7�e�@nQ���}��)�l:��*���J�9��>:�)c�A�I��PHF뒥�f|%��A=c��Ti��Q_Zs��Uϙ�/H����.�r{��h�1�3��������7#�r��E��G03\bKDM�v�?������Y�gpD?O�Zv�P���+�?5:K��F�\*t1��5gS�De�<�����\��,�����^��ɚl�4kQ��듄V"����#�1��l���^��M-�	�q-�ҏm�H�7C~
�����X�h��)/��N6�V�7�������[��>.UøhA�ӽ�#m�A����L��7j�wf.$��Z9̿�`�����VfD)�bA8��B�J</��e�6��V�7�u��՝/X�܀�Ra^CTK�9���|v�)���U������&���ֿ5�ěj�]��� AMܱ*P�{��� �*���,�N�q�q%x|��R?����M8��$]<[>!(T�ZC~)��!�Sy���,Ǟ<۠�&,�{��O����?,4��^�S��2�32��%
�[#�ﾱ�)��
!���Lt�0�
���aJ�(�2�W���y��8Q���^#���<�|B�mð�ۇ�s䃸��xv
�˂<���4<�U32��'��c�7?ME���f��P�`R�����p��Y�q��~af���nQYZ��6�6J� 5R� ���Aj{:E���������)����)<�� ���qC���_>�8��x ����ތL�V�`�#���M�4��;�L*��'�°�-J#%��/�ق�'����VP�դdo�d1�P�0\������o�ܸ��.[}��"���п�%V�W���u-YyM���D$��D��������O����e@��6n>��S��l���9pt�vQφ�<�IF�����ֶ���]�.��������~e��#�yLdrq��xI�J(�� ��������'���/N!�Crb��/������G��d�X�6Z)�n��s��H����?�3\����Ʌ��5�/�XخZ*ܨ������J�:=k�P�-��1��G|D����jm�$@�+�f>�!	8�#�Q�l�����Nlǃ��X��!P�/J��E���^7�N)~�-4�"6��.3���!1�?�ep���Д3��p���~T����
`֦&H�"ץ��1��ּ믓4�{�<d.2qË��Z��;�`;��t�_��%a�NV��u����"_ຨ^*���W�#k�ı�Ar��-�j�9� �[�p ^?s���o���gh���N�0�z)�P���������aX�b���_��U�=_c���[��c��F�a�/zK�f�9��o}l!�c"_&"I�,�m��V������j\;4��P`㜖�sA��2��4�R����.L	�� �ō��&`w5A�G��V�:�2��G��S0�|Ҽ��o��-^�n"�7M]�^����p����)��N���r��P�&���R7��8)3�OU�n�� ��wI-�l��@E���9�����y�O��+!F� ��@�����VJ:�q��	�V�g��#���Gz;�LR�,=e_y�/��/	�~��_ݜ��b�휪P*�B�0?��{2j�JU�Ny�!�=�T:.��6�g|�T�4����\Ѓ����I��԰/	b���NR�4��\nc4LN��L_�M�}�����.����Z��^߅hsެ�����H��nB8�l�K���H��Im@��Piت	���Pyq����VMa�T������K��i�Z�i�H��w��OJ��9��������m?�����,hfĐ�.,�p� ��I�Z�w�A�g9�K>y�4R�W�\T�lTS2�3C�c;};��v�&��`Y��-?��������R^}���r<��e���p
X_�F�k��i�?Zǎ.�	��S����4���9F�,!�����'击p"��O2��ZBv�H�85�{�i�h�86)z�����jq|WP�b��ͳJ"��;�?�@C�Kmw*�q�����`�9҃�-��FZr�#����S�Jl�W-#��o�5�jD+��̲%e�! ��٧���N���C�!_�bU_q��6�k8�qa^I(r��A`6�<&���9L��A�
p�{6Y't��u�,��h�v��˔�B�=��!�h���tQ��z=3�w��c�)׀��������
x{�~�9H9��*��3=<L���,zf�E�`�/�����Q�x�b�`�^U��d��[f�ɗp��\�����ZS���ޢ� �[Q/��i �OkW�B�F�z��U���	pL*j�M��4��|%N�{���̚z^�%2�&څs'n�4�N����n=���Y����K�mmxq�j�^�$o^��cs	�������Fג�\�Cx��`d0�Z��%pq�6ftiq;�C}c6�F����ۥA�L�������ţR�S��
i�R\X��v��'����Ye��>��mU� H'W��X��=�Ғ`6����