XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���uS"�ӳ���H<(�c����l>/=�'A�ݪ��R:5�u0��Z�Y��( _׳�b�U��~�t�w�}���v�?�Y�qY>���mV~��0q�΃�C�ai�`7x�����:��`�8�t�̀Ǔ|�j8|�g���݁@M�u;���Sh�I�K��6�p�o$0��1�aD'\�-�T�jsz�B �Zc�����E��%qS�W�2Ʌc&G�YI2��Tpl�,�a4?����*J�KGKcQJ��.��*N�~Og�+�{Œu2��BdO���+�������W���w�'�t�U�7��
Z�W4m0�S��l�Q��B�t��A� \���S�Y�fM՜�YzX��K-@��d��7vԀV�ܓ�]��Ţ��r'>�SzJp�w��q)�߆�*��Qe�;���t3#���:�؟�Jz�'6�7�.�YT���$��#�igkT�p�2�����=>[Ԡʄj'yVAg�9|������W��%�0�_�[�P`n�6�_��
����~1�c;џi�k�n�v����_�͉�Gg��(���f�-�Ȣt�����~�H�Z��V��?2�w��/Nj毃����7Ũ����cj�:?�]w �J��������*!F+`�6��Ѐ8W��7&B�9�Ҕ}�Lt�H�:Kp]iʭ
�o��k�z{k���;�����Hj��m�#ܚ/���tٰ����T~�u̩�/R����"S��?���$�·\XlxVHYEB    fa00    2620�5��r��3�!�6���&��]j����j�q��a�+{�P����0Y%�&5��~f��mF!c�$�s3�QV!om���Hk�p�cp�՞n�Mޜ��jʎd{t`4nWt-���&yRr�2EU�N {��d���l]�\?�.9[Ũ�tk�{.D?�Z���AQ�o� ټr���,��hߧ�p�@�J���{0��Ϝ}���	�������E��;M�ݗ'�cM��ɍ���Q��e^>+� �laJ���_�e���% |n���Ȩ!�c����E �j�x9F�~��%�އ�S�=��?I���
����9zpU�-$����(X"Ư�l��as���%m�)]y�+��1�����`vc��A��'����/Uuk0бh����� �`%T�A�5t^p�y(Z�iDq$�雍�&��#�g3�
��p����^�D;p�:3�5��jVy��J}RPi��^����z[���8yN���>�>W�n���d|m�y��F�}�X���/�Q;1�m��a�k��XR�Tnu��SސX�"PH80]·�<�vep�[@�['Vc��0_)�/g)��ǀrs��ٺK!4_����7`,���eM[��2�'Z/�������}���]ȡ�ۀnI'�E���&vp�<�s�N�˅�j5ԁ�EA��t[����'3��9����֕U|��B�
�ԭ�A���:z}�����Ei���5�R�<5@�Y�qU�f�%h)�y����k���xq�����BL��\��?�0y��`��R�ga�VK���\�R:QȆ��<��p*�	s�&;�~�?#��K���_�un��z%��.��FR.�X"�p���sY�}�;N��,h!���&��>M�c7ﭾ&�z���\�]D��qt���6QN�kOv׽$����r~DJ�3z�����q �<ͯ��֜#+�%���L4P�"f���e�zdC�P-����4����"_A� �2��l<A��xt��<�x%�����
0�˴0���a�Y�Z�rO}������;��T#�^
�[���i.�T�w�O�o#$�E�P�(<-1��ɜ|7��
��������\��h��vhr������Ej��ZAHZ�/q����v.";�1/�f��8�V�U�:h�0&�aZ���M�@N������&�p��HZC8]0��&3���n�c�������6_[��̄~�@���gu�N�L�^ۊ�?�9q�b�>�K������Tj�E�{��RWJ���\Ѡ-O����r��
����Y�t��9�Q���������"XZ�f���"%HS{���M����';s��\��j�c�����R�*ʞ%����8�\��Щ�����X��rB��������\L�Β~�a�)�;��������\�ra���ѣ�r.��p�M�Fd4ѽ}k�17K���ɉ��(�2�y������zԦ��}�}�.�ZX�?u/�J�Y�C�����&��֣h�5a�oN>lъ����Bs�o5���K�,����XW���ҫ&�� �؟L�����yU��i��w)_p7[h�pv�K�a�j��s.���P�[�<�E�ݱ1m�Y�ሽa����C����N������R��C1�R�q������՝��%'�n>i�:�:܈Ҩ��qU�O��Wz8;�;L���w��/S�hŝt�g4�R�\U�l~j�yX�-�"i��rӎ�r/_�Ɇ!�9�G�͔��}��O����Y�]*��Hs���{$ۣ�]�K�����������8�o�4����L��,�"��v��T�V���b7e�͛%ml��4|b���Ғ�866�ވ�${J�{��dCi"Z�� ^G�²ZDB�N��'�]J�1��H�δ\�;�Q7Ԝ@�D�/2��C3ɧi�t�"B�d'���ca�i�Tl_�y	��u�cJ�&�0p)!^|jܾ	����Ȼ��te����
z�={�|��O�����V�����iw���bf�(�D�W�@����PT
��X��4?��u��E,ĕpiQS��-�epĽSl��H�go��Q��P�MA���GSƥgpu|��I8x���3��������������[��c��)� �u�X�e� د�������='�E]͌��f�$�h�����o�[���0�Ɛ���rF�9dy"�4�zf�C/��6��3���E��Po�\�*a{��]�E�� &
c�/D �� �l\E:M�J����,�4�q��N�?0�8'e�ɇ�M�`.�s%�pHo��M��f�5V���Gҥ��N�� � �!dRX��Kީb|%���#��L�&Q%,��ߴ����O�,�[	��m$��QJ{P1$��_&�F����|Po�]Ŧ�f���'?h=�E�lm�p��oĮ�Wf<��݃eݶ��<�:C��oy�4�x�����ΐT�#��gV�}h�� �����bn�
IS�xQ`}Ae(�ӽ�?����6#ׅÊ���h�`��I��W�Ө�6n�d��e,	����E�|�v.`��D����G֏d,�m����5�]��3�@�ђ� =w`\ �V�;z-�=�����ې)�LO���Q��[W���}p�@ȵ���K�`�Xl�-�=�3�{@|`��]���)o!�`�<�V���~q�u� �(�~L	��U�ī�,�؀�M:������kX�x�G�~��moL��Lv�1]�Z�B �|d���Q��f慘�ɨ�׮.1��FI��,g[G��+�?C�/=�R}$�=o̆	c�וS��<��L	�O�3�$/G�d�P�g�g�4�dB]�G�t�k',���KΫ�>�� �F�F�If�{s�fM[�ƿc�d9|U�LM���������F��Na(��\�l��H�ڧ��+��t��4ƸiK � �f�!]|`!3s������AK�AxH�������"�U@f���	f;�~�<����u�G_.%X뒞�b!汏x���Q�'�V��,(�ׇ%S��+��K�P=7?*|e�������/(.��>g�k��Ώ1&�zF#=���T����3qS⛌l��U~+��n$����Z�LFX��]+���X�G�5C378�S�=����
y�er���+	�8���o�Fw{t]�"�����RZ���� ���we�����,�X1�38��j����_��Iʶ�O��k�i#6	�uG�̯K���;n%t\�ۢ���%1�R��8H+����eԑϿ$����^��5�QH��(�u��#O'`�L�V*/���y��Y��Ch�D�z[=�Szt��:#_W��S	��A�S��7��N�������	�FN�o(X�Fq���x(0�{�q�	�m0D�4�*�h��68!���a�/��r���rR�7Gu���.E��ل������z_Ìv�pt�h�p�j�Q������Hl��0���Y\Y�D	������35`�,��O��cǯߪԪ�Ӽ�E�3�}�t�C ����i��'��DT|�o�HX��st��Q��j�/�t��/7,S��<�����;���xQ^Շ`ܜӂ��s.��z�,?�m *��x�8�j�Ksx���I���KP��\��㭇r�FKo4�"%�5�^Y�r�S��.�^Ѽ��ݜ�-%q�����&9@� C�1i9���~�J/ۂ��!�1BS��i��[x�`�D�t��pqV�>�3w|\+W;$��[��㛟��;N�<�|M���m&��Pc7S@Q�QD�+<
Q2�a}�h:�>9b��`q<��d�"X���@q��9C�˳�yz7�ќ�w&t�Y�������Ht7�����S2���Ms�=˖��8�mKx��Ϟp�b1o�ĬZ�p̴��4�ջ��Ĳ=?��D0_��s1+L���!Q��Ab7���_��sd�uZ8�߬l��_֡+6|`�k@p٧#�儦�� �T\G1�?+�u�x�C�w3�|m����w�w���d֋������/�My4�eMГ�/�����9,�ܪ0����n/;�n�HO����u��S�/��ˠ#�2��O�7� �g!o�Z��8� �(��0.�qA28ѡ ^�4\3pY��76��V?B&�Ž��ȼZ�x�˘��y�mѳg޾�s�D`܎������&d����ې�o�/]�v^*<�Y[Ƹz�Da=�G��#�m�褐*B�� /�(
l�74)��o��/���V��)�0�
G�F��L]r�_S�݌7�v��_�!�L�i�HH?J�BQ�CNw�/+�2�h�G��D�����U���.��]GeG��v/�����v�9)�c\�R�8�n��/���=��n������ �_q)�n��8Y��]c�G�'Q6���`2�v~Ν��_��H����CPx<�
�#�}�*��rCI����%a��@�~/��_2�����x��uӪ	��
�C1�*cQQ�KT+(�饢���3��G||�'^I�.�}��r'��em� ������o3k�%��"�J�o�<,E[h��"��w�ѿ�k��	T��Z�3��W�(u8O������Qz�T�̻ڞ��CƂ}����{�Q%�3jG�ߞ��!;q˘����׆�{�bi���*�v��<���FQ��]���ǯi輠\Ƚ��v� ~�E���)H���H���4*��
}��3n��0��d0���2�0{�v��#�E��O�=gwW�/� ung���	���kDc��J�򪰁1M�-�|k�������ދ6s�T8�6�e�	;DȒ?�UYg���Nu������C�����W~�v�Z�s��/^��)���b՛�ؽ�)'d-�y	��jg
���e��>/����[Bj�����7�!(���mV��JN�h���w�K`���c�����>�`��'i$��rH�݄s��';�sC�AH�c�D�%]䥺���s����z^o�b��6i���W
���ȹt2>��6�7V��,�_9-����]9����L���ح��ק�B��	e,�QC���{%֚�,��<�>#~M�u�>>�J�����t��ƥ6��(CD_6�=�kzr���Cv�G���$��� ���Gt����Fv%��5`h�f�1FU/d����b�T6�C>ŵ�P̷cE�� ����֐�^�La�E�v8��jW`�0��E��$�o���L�-c�É'��� L6��7�b�w��V���fd�;��ߝ�F�к�����F�������{P7F8~�Ѝ��$#�A��fo�:>֊�k�YA�)+�HrX] ��@f�gkUb�̗	��U�>�7��2�� ���&�n����i_����}�8�����/u�?T\�c�i��ڏx,A2-�9�YF>����Bbr4
�yš��/�����(4�QV��>ި�x� .��A`WQT�X�g�3��S��.-w�ֲ�(ڲ�lV�O駭��8���W���=fs�R�֒Q��8�Sq�C���&6r�D�=D��ߔb���W�c��cW6��������Ը��oE}~s��{���c~����J�/2�m?/��Dl)��WWA	�W�he7��X�}�r��gNi��@>@�[��[��i��{�>��w@4�{`^ޞvI�N�	m�(��y���WY4�|���K��4�Ac�*Y�� �<�٬0�c�t�=�]n*���d�`�h
|��cɇ�x��\��U#~���Mzn���B�n������rPvr��C~K��;�������w�]���$d��8���w*�/g�c	K�)��ښ��$��'b��_����6h�{��x�aMua���Ta�k�pIJ�Sb�����q��!��~d�M��L�_�2����	^8�<��8��T�L�^T���?��u~�ІGHb��W.��)�.�����9�N {h�w�/��F�UY�S��<�!;;�\��e6*�š��jeX����F4�?J�؊=t���d�Y��1ң��d�ه&�p-���ܘ��E���<�m��梬�}���GDӡƷ+�W�)K��dҖ��W���Vq"ؖ��Ch��aw��f〵_�~�C����I�H�dy4Y�=a���ja~�t�4t=b&�1ͣ��3��y*�;Y�F!��|DBbt�4�EA�k�"KT?�e5<��f�:�����w¾U�Ǽ;i�_`/l�~�G�y�-���A[(��{�0��j0^��c2 �Rړ�m���H8_:�� ��z�o���<*&�q�}& �ߛ���lP�mw>�C����K����Q��a%WW����o%Ӟ�0��4��w��P�Y�%Iu�ZT��E��O����G;EF��Zf�Ok��#<|7^��	�h��?�k��KN�����v�V�R��x�t�=f�u,��O���"��⠯���k��+��7�����|�L�3��\)�t������"=w��T@��H�k���,��9{��ԄW�#��ܿx�߃��j:KkX��&h���V�=�G}sOfRusGp�I�g��B���iVa���٭&̵�6��P� ��z>]���Z�i���6՜)3�x�O����U˴��comQX��M]�؄
�g��=�:�����鄖;g����0�L[��/;Z��,���������<T����)�m16������i�m�_Z;#܏��t����h��v�Y��H$�i�IX�}���A�QR��y2���Ba���Y�+�)�NtH�����U]�sIC����v�K��B�"��4���`͠WN��3Cd�:��#�ۚ:
j��y�%q���D1�j�b�Gg����5�<9���*^�β���#��y~�qR�{`gn�F}��K(�*ׯt^�T>��	�Եu.@<QA�!<�Ϸ���C8��-�}q�~��'��e6�T��/W�'�vU��qP?��yE��'ߓ�ze��,�Sԡ�"j�#�B����?)O�K�J�M�u>x]�P�ş�[\yƏzE��!ڃ��j��������)���;dD;? h�A��q�%�$e�e>�xA�}�d�[�JK��I󄖡�;��u���ZY`�l�Rf7��~!~"��m Yն9zI�n�� �H$�;�S'QuV�C�g��W�=�E=*�s$�}�Dt!�F�k��@�@���Dxz���;�r�|�z��Z
AEO���;lm麕��Z'�����&)���1�T�צ�cqDzg����R��$��eV�L�������sv5�!T��f;\N6>>��ޭ>��FfL���Wm�(J<q8�٥��{;�';c<��Xx-�]��0�3-�8�����c�E/{�q�0��{�Tܗչ ���8��1�!ߑY�N�_��tאx��ئ�흉�Ӽ�;�LY;XY�j9�/�˶<�6�
L$a<�>E�A6��8
9?���1n��k&L�Q�\�� هɸ���hX[ʁ�A�f���ց�mL�4���%XLʃ��\-�#�3��W\�3<�9��X�NN�S$bw�W"ã��*[;5����>#"{�c���?5L���a�$H��D��P�Әҙҽ.������hfB�ꩱ�Z6�lZb�V��Uj�Dr�-Ex��W:�hRg<t�m>R��b-6��:͚�8k�^��*s�ڋ3�����S���i��n��S�s���ƪ�,Iy���:3��o��lUSv"AX�e�������exQn۽Y)������{�u��ln{Z���xU�3�<��P�����6���$1���L� ���P�'�"D�F�ta'��}�Hu]�S%��h"�AC�8
aԯl-�`�������lG�q�7�}�����!��K3�����B�Ag_��W��M�J���%�8�s+��ŭa(�qFY�԰:Uh�0��|~X���u�ku �[t�,��C�aV$�d���>+r��_�g���J�V��t{�)�L�B�)�sz�W�g���͍L�s��ĝ��G�MU�Z�N)�D:JOB6`}q+̔;c��S~�?�����7�5Ba��m�~N�7f� '������*�
�΂FK��&*d{�'Q���fU$\���~���'�b]�w��I,����G���}�గ�J<�1��jR����{�����/�/��[�nB���6}#��uSVs6,��E��l{9��i�����dZoW� ���>��*!���<���|�#�d���P٦�*�6/�Ȝ)�C�F�JAо���ڲ.�aә\�;ner���	��DI��S�4VJ��"�H<!�����ri�H�Wm(
�:���r�TbI��{?����Ґ�a[��m8O[3���g��`�u"��DD,�I}]^7�}����5<
�v�^�����9��J�<U5ũ�@���3�e(�xt���{L�@�77
O���o�P����Y�:х�����5�!�po�et�LxT�_:�zsaǿM�f�u6� %!�	*��������Ք�_ā���6��'z/Ƞ��
�f���V�iA"�+�gT:�h��&&t���T��9T����])�����\ޠ�!4��F�ٶLn6���-�E���J�A���fR�i���\O����Kc[SY���"��6�ٴ�G�N�{����M�s�����6>=�_4�7�}~7\����t�?l���ʼ�퉿�����MYk�#J�ߌ�t�7����;��7�H�	�w��Ar�V;i��,�|�]��2i�9��޵O�mƹ���n�_����Z߀�o��9�m�=���"]��N�����,7Bw��1u\�IG�|�kP�)��p(m����C����1�7Ԙ�45M�`��XND-���[��d�) �*��~]+J(��O��'x8P��z'�����Qu��*R2\0��v��<"��62�CD��)�A��S_�����xrx��փ�r�o�Xs@ƨd{��p��7/�7KPw�rr���'X6����}tf��44���N���"?����V#�q
m�%i�	�������Ba�;�N�FjW%���Y�b���4"
FU�O�؄���٪h{r7N[_�xד��8Vt��}G��uq$�!1���?��	&�)C��3��^�/h������s]|y�uu��{qS�-��0h)�䖒�=ڹ�p��
!��Ao���Н>Fz�߆�I�9�03�c�u O+��C)��"3�k:�K��D���W��z
�S��\�ɣ�nG
W� Y�̌��*$��㼑v�E�|Y3���$�L���Dk� ��y�<�v*�5�Aq��E�{U��c7�N�` ط��g��k{�1�Ӳ�|���6�xJ��r/���`\�#�|Y�2HpL����=A�N��q' ��ќmQ%�h�a��=����R�]��ȥS�r[Bn�8lz�e@�z]Ao�D�� 625�C�{^�i�N�+��A��}�i�+̂���<5])�C�Ԇ�����_����.�'�¡
���G!u��akB14k��'w�ު��_�Xax���Υ�����FU8�XlxVHYEB    37e1     ba0>"~�����7�~l1��w�� �ێ��:�Y�ܾ�{Ҵ4}mMshS��y�~�azᕝ�F�����E�J��a$��MT7&���1:y��,oy�~F��9W0��c���>-��v��Ͷ�{��i���3r�7�hq����:�5	����f.G��a
�r����{�"'��`(�%X�<֝�5��`����*x��Ջcz�~'Ձl���Ǉ_J''i�
w���C`�tWP.�J_��&=��E#K�'!Ղ_p�����ǝA	O��o��-{ٕe�BF��6xf���:��A��~������4+yz��������"�l	��ٮ}�Һ�Ѿ.����4!������'Puw����o;�1`���������3��$��*um��m�����WlZL��Z�	M�g�毀kI�N☝l�����r��"Ҋ[��Z.~�v�h�:��w���s��O�ۃ �����ݯf���*M7�P+�M�����׊�r�Ć'�y^/*�W�����2ф�V�c�a�I� 6�5����3*�x�sNFyt.9�/U �Ό�����4f�njlD%�*�&�I�q���]��������$]���;~�l�J��A��]If$�L�W#4lt>|�x+�Բl��
ir�j��Yˀ;��t�"���*}����s���o��ޒmHM��*3���f����Ō���vG��
��y��2���E���G3t �ǆh�z���m�Jh�L��u��L��H��<�̉��IJ]a���̆������}��[�&\b^N}}�����JJ�2٫�=�6����\�s/��<�,�;��[)R�64�$�i:	7�F�ݛ���]�ޔ����e�����%;� ������s N�7���#oe���SAI���>[��7�B[���y,�972l�����M�{(�"�	w�5���!S�}�Jo3JU�A� lw�G]p�c4�a|�ڋwj��[�bI0�h�}�7��{Y0`�sl���M�A����i���[�\��lB$��c*�=�8��5%�'���t�GR�Ŷ"�t�/⬾����2p�#�C�o ��ܲ�����>BQZ��(2@�I|_���H��U�L��վ@�sm�2@�A*�)c�HlO���H��:(�Bib8����-e��R�EU�z� ��p�����}����C�8;�W�œd�����͐����S��NkF�<Y�	���28�����g��7��#�0��\���kf�a0p>�6ܸ-Tg�%�s	�/C���c�! 	��v`�:j=��}as戾�<.��.��f�L�!l��h�?S,�~��R�����-��sAS/3�+�� 4I>hхW��76�p�ߕE�lp��>KE����Ĉ�A=��Io����V7��9`�P�i�/���:� L5�{��E��`�&K(�"��auA�E,�.G�4![;���2���k'6�h�g��*i?y�~\�>� a��ub^�J�<i{����ܟR�wz(UW�'�K(�u�i��B���Ĉ�X�E�
~�@�;N��y�%��5|2~Rz�t`�Q��8��8��'��<=FP�zӿ&�/ϸs�Qkp�>?1�VL��*��-!���p�X�/΅�ye��כ�i��$��8f�wn�������~�)�x6�9�[�
s<݄�4�,W�"+Oͪ������\�ܿG6bQ�+��x3O�KE��k��F]ȵy��/af�_A�<H�I�QW̑��O_���">��[D/|3�}ˣ�K|6(�'������W7�[�`�p4�k�]������N�<����[�UD� �\s<ay�Q$&�[���J7�f�l�q�{���=�;�+���z�@�v�=!�I$���c`�!X���c����w�	^k�X��U��<�<�r�V���my����N��j���:�5C���Smd��^������ �yL��I�zw[ƿ��N�+��m� T4V�*g���5��b���M���g�-�U�|�[�E�/v�R�� bԁݍ4�[m���}N���h���F8PxD���~��p����B":�55�}�$*~�+>��h��O�d��gM��c9��l�E�\�q�wm=oQ��~��k0Dy�y�g��l���l���	���o�@���}f���f���Z�r�=�K;��.{YG�:���d����p������2���ƙr�ڂ��Y&4ma6�u�����=�9w��n��*.t��-�K��H�4_6������̬O����)O~5R"'b!��穏*D��^��U}o����D[��H�5Πܥ���a+_����m"&H�~�p�K��ln��Bm��y&�9���y��*ޤ����6%FD��o��VH'���'��C�vv��?�,_BZ S;�%��Xg���64;?tRI�ʅ����	��x��}?*`���vO�m5;���c��#X�E;�����a�S���]�h����9%�A�Jrla<�¨�;7�V�R+�-���K���[N���;@S�P�o��#ǙR���cu9����)e�ᅡ��H���4P|8�a�K*�G�n{%�(����;�̎�^�S�w�����,���	d2�^��h���wԪcih��#��|L�*n���ҿp?疂$�+�y��d%֓��dp���(6>��E�YB������߇@�D&���へ��Z�bs���Ҙ�2amf�P���Qݯ9#!��d�m��E�ѡP	������͊�/T�����l.�z^b�O�R�~+���n@W�͖�ܖȜ�d�\<�t���q���Q�wj8�>>қ�	����k�xv�.����WN/���vj�;>?�\�S\��(i�V�﬽�`��7!B�G�8�W"Jy�x�p�׉r