XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4珀�w��F���^5�R�	����������r`o�U�5�����r��	��6�Zlȼ�:ڒc� �ps�����e��<T	aH5����d^A^r)R��\�Ŋ�.z9M�íʠ-��J(?hq1�|n��~_,��9��ыa���I�����	�
�������<ۜ��/2p�G�J%ü��@�u��=i߼~DYtn5s��Y3J&Ƴ��q�p�jt�	U���l�?���y8fJ��![�|��d�1�X�P�T�pI��<jl51׼!%p%�/J;��Ե:�	�(7�T���F��b_�^^��|��ȶ��$���Ҩ�5����~�cl6����"dx�}ӭ�?ޥ
ؗk?y�|�n�$�����u2ĽQuj�X�Ӂ0�K��?���y���oI�A
.p��	F�M����,Ao�G�� ����"j���Q��ڷ�� �(� hC��,SO�r�J�Q�)�Q��g�sV
�L�H���_ʷ������E��d
)��uٰr�c���,Dڕt��c��Vg��Qiz"�
��۬���?O�$�M��ǂ���a��\�`�V~+�0M*��d�ژ~)4ZC�ag��$�Wq��������� ��EJO���gI;���S��N�2�k���`o��4h�}�z�9]t
O��W�sP�����9�ɼK���Ϊ�b��v)�nQ��{:5`�����[(AG���&lR�`��0��sq�ld��V
@��"���2U<�a7(ݙ���@RT��ȒXlxVHYEB    203f     a60��!\����4���k!WϮ_��j.�d9[AS��R��Ȍ�f%�ɯ0���"�x������\�vO��,����pL��|F��/�{3�P��X5�9���4���W�^&c׊�(k��`c�&��pX:z����`�%�0����I|�$N�_no�a�tI��m�?:��)��Yy�z�΂P_����,��#pT{k��CSS��I6o*,:��������e~�L�����Q y�U����Y'u�ZJX�|g��|�O7��)&[i�sdd
ӿ�%U�T����:���U;G6��c��Q3&q���⹞V��w+��6%��I�"��56K
���G"M���4!��&G��neq��<�\�6~��oŶ�/ߎ Tw~w�}�=+��Q'gB4X��^��7S�/z��s Mv���1�5z��H���ح=����8���h̩���<�y
f���F��<D�$����|���|����M��+���dv[�I���J߅{���p��݈��)P�x�ڏ��z �T:������Xb���!#"�id-M���Bh��?���<�}3�{���Y�y^KP�9,��N)e�P�D�<�1h 2�k�����bۖ��;i�[C���������ü�D�F
��{�����y��e���=�ҽ|�A�z! \�G'�f��93x8�65��ůVK��ݒY�o��F�®����e�Cح������`\����M�ԍ��S���.�@�5F�6���ĉ^J��������T�MbHe?6�)�ʔ\��Ĩp+>�l��UNZ��ٞz���|�P��!UW
ܽdwph
�~LhJ�OJ�8%�'(���>�2mM��W��U��D���6<g�M�&�&W����=fae�,"Gc"	���(��	�s"���0(M!;����Ǎ���2/#뻐�/0qm�ުh̗��]�ҵ6���*�*�*��/��@c���	R�ð���&���#�}){���3��Xgڢ�M��-��Tf7�A�Խ��p����3F21�ǳ���*�e: �Κ�;�C:m�G�xX��E,�j�샎�
�ށ�u�̛�L�E��v YJ�Q�q'��&D*�By�r0�ռŚw�p+YƩ{�%.#�#�u~#9�W)DM>C����4(��z�pE��VO���8��Qb��c��J�fҡA�hnd���jm�q?)`*A=�X:]I�Rx�
r ��&lP�5h�N1���o�x�p����&L{Q�IP�>u�sae+N�*�����Z��E�����X4�k�T�FEp� Wi$&�q���O���&�����c�����6i�uv%�o]�
��r�[�s������9��0�6ذ*�ǋ^j�hU����pگ����� �}P��)��Q�=D=ɞ���b�k���Z���[HQ^�l���g����AѨ���8�P�bY��^R�i��f�2'`y�[Hx�Wo��<B)�b��.3��fF�~]�^��Mģmb2?� �� t�+��f�!�^��x��I���8�y �4P�����W�������vl�����[>z(�4UĈ�Ԉj��,<�I�������,���7��L�+��}.�1������`rC;���],+7^{���i�A�xI��+��x��� ˞�&��4����n�-ٮ�)Sa��YxD�۫f�R@�q���	���E�%Q-�<L}"@)���Le���������@�:u/�*疆漨X���O){�x
;;��S��Ϛw�r���"�����G��p	5���L57_����� k���Z,L}޺);r�%4L���>ڶ�9��6�� �>oI,�8}7�˲y^��q�c�l�Y-\J*\��3;�/�y�H��J��d =P�\	�Ev��9��������"��I6?�Š )���bYu"V�j�> X�vs�a�D�6��g�7�k�E>�l�����/�.�,���B�-��k�@VYa���&#�(��Ibȡ_���kA�l�5m�/{��r�=�le&py�S|���N�@B�LD�]LD��0����Rw]P$�<��tF�Z/��̌^MM?K�w���tQ@����3�kE�r͡|�LP�n6�h:˔S��W�(�I�w��b�2/��
�a6rx�ވ�Pʪ�#���Qw~ѝ�'7a�6!��Qʢ}�~�U�� ��U�@w+��?�	'-P ,\AgV��N��{�j
�Qݣ0j�N�
,A�E7A�TiP�Z��t��#��pSh0�?R,RE>'��T�u߶~D$��2,������N(���-�8��+�,�q��j�DH���Lk�'��*e�$S����J�@�Q�+b;�g�8�r�ld�bۜs�l5�]����[72�><�|�/��<Zش��C�Hֹ�b�ü~8�zA��vNÓ;�~�Yi����32Aat��9=�~��]H��f3��3�T+�ᚌ��`αf�i���i�UA��<�_sY�#v���ν�|���g�'��4(��hR<����$�-%��	�y� ����_i{8p��b�k��驲k�*���:�P'���Sf�9�G4h�����U:���Y�?�����A�`��0��@�M�E�/`����W,5