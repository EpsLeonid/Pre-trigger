XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r#�tf�y��i[�:A�덉Q|��L@���KT �%�
�1�k�IEc����I�	��i�Xvq;vevR�$;5A���,x���6��V�k�ھ~qaOͨ����$�[���A����� ]n��,��<�l�. J��UJJVo/������}��9+�����d�";���c�Y���ܾ�N�=���i��D�s�0�x!7�O���Q��X�X�=��_� ��C���϶���a���"��=�:�K%c���"��O_:�w����y�>>+����ꋯ�����?(̚�B*s�i�M	�c:��_/�f���	���LQ;
n��"���M�:�!&R�'�����մ<���r� �w;%��Wd'4�'�e�n�:�	E�$8�b��=V^y�/ ��Zi �ePG��y"����\�(���R��$ĺ�9v��:[���R�4y��o�,�Z�V�D�U��&\W[��i�kVpRO�!�L98oP�R�"�  �?="C�����]1���R_wb,O_���n�WF��*Ӟ�.Q����v#��:� ߐ��΄�Ǘ���3���K~�u����[���N, �8�g�?��"�8�,ܿu����S<r�hb��"v�6�
^I�O�Q|1��iwm��.%r�H���MNw���e�
H"�����r����o�dFEB5��>پ��������Ҷ����Tc�0MVml
_!ߢ
��RU2����N�mE�f�yZg[���@f'�WXlxVHYEB    47d6    1030zcC�B-�Q���4!�j�[��!�v%�[������8��٤{��}jd�{���?;��(Ӏ:��2��<���{s��t�7�<R�� ���q6�V��! )��ZR����8���sH\��ݮ��:���֟���:Qdw����$ѕ\���C�znRմ��0���ڰ��n&`�fx8��0%����9�a�C�>+ꨮT� �9����)��d�#��5�?�p�s�#����j�83�*�O4�Q�W��E5,��nVRz�����8;+���*ŻX#$�)ʉ=�4��b��Kb5��������a��s_P�c�mV8ZaV+�@0���Hz�T����O��O����^]ގ���{�u��^ �|ź{�ZI����c��=H"�i;n&��Z%��?~h�>�Kd�ՙ����
и�Ɓ��\���_B�4ؐ�mN�K/�k ZP�7�٭��.k\��Y���Y�J;�����X�(��i��\�-:�zw\��,�1|n�=�����8�ű8���=R䠻�q��II�<���H��zEU��(��^�WD���F�&���g��B�H��>�����8����x�`$���F��頍WB�#'ُ�<L�e=�t���C��t�T��-/���ۻMhX���p�������3�
�� S^N�g���*aL�,�B1�o���@��y@(8�2���#�A�-G��_N>�Fӭ���'�#=�~�kC\����u;��8/�譄��&vW\0�!o��s�#�z����n�|?�9��='/�3'dc/Gv4�"��;��T���"X�b49�R�D���)(N#J��-E�}��b18�=~�o=�'��/DX��#�nEg��sz�SZhķ�7�t�?��ʵ�`���2U��`4K�f_/��ڇ�Y��,f�<ڛ���J<_ʍ�_/�����)]���<�.��nƾ엍���\���o]?ؘA\\�wG`|��"���
�/���[�-� �r� u6������#��5��o�����ř��69�c�̢��GN�#Dӊ.���pC}r�R���͑n,Wz� *1�12�����U���(������#���Q�[�������7~#�QL�l��7��Y�������K�_keO�i�����C�X,qL(��3t�����Pf�3%����ՒT�ٳ���(���!2H:%ÆOV��c�ԋ�A�{s�Ż��wA���Fkв�����+���nk�����G:�h�ШRxƦ8Hm�Y�u��B 8��ǃ��m s,���6�?��vyӢ'�R��Sf�qE��Y���I�{K��*j�:��.͌�ʳ#��@���6���X��m�L_4��jS a���c�R��N��K�ѥ��F��vn�  �I�W_Z�4��D�|�?QMY��OȈ���׃��-��39v+�#����sp�UNlfճG�moD)���L�HP�h�()[1�-/	��rDG��d]!TUW��m�12Ƞ�PH`��t��_�����3}�f��@v��S]��@���fZzr^S�b�]RX��}t 	U���p���iL�s� M�D�����H��NA/n�D�S6Mbg�˃Ƽ��b[5xԞKS�Rw�ϰo^H��U� ů��}����U��jc���!��Cu#u5�hX8��O�>�h/6O�s&�!�t\����"�L�>�KQ6-��iL�Ņ����~-.4;N�`�E�>
����<�X,ϓ2���b�1
�aG �]�S�X����+3pe*���U���n5��u*����*����2u�*�t<��z)f��4}R������>�����"�g/��Y�r�9�����_fMY���ݭG>�w�1�e����W�(7��4�pt���v�rD��#G��I�S��1ATf$��4>��G���H�
L�5��<L>�`t�� ^��d<(�?���&�sQxXp �Z�X6�03K��?�ib�00%�m�G��ͥQ�u�N��צ���Ռ�d�T ��|��FM�}���Dv�-ʮ�%���-��Yj[�<u�����F2��շ	Iک�h�������c��d�"����X�y��.8��=H����u�,\�r�	��S�_޸�1�=������F�.ଇ]�w�(n|㜽o�W�n҉D�ݕ!����B���6���@Kd�����en��Z�bX�B�<� �6�j�>�?������=��72�e)���^�,�/�fɈ:�}<ߒg���;��x�v�D�?�B�h��޸ߍ��嫹2���ꈚ0ǧ�_G*�ap�P�JP���w���6�����i��^�!��9&<��g��F��I2)o�7	u_�Dt��9�.@6�ߺ��K`�	m���z�^��C��Ϲ�<�f�7l������H$D.�tԹ�>�l��rI�/0S�+ͷL&�<�t�*�����`/Q��/�8A.Bp����kG����T���j�O_���\Z-	�[>?o�㞾%&�V�	�y]m!��)��I�I��a�d0��@JY�e����O��j�Vx�]?މ���"Uح�	��f׀�����v-8��Ǭ��|֛ڑa��������$��♢H2�DH�E��ɬ�F�W���_�Cv�VAc�R����r�m0�p�m�1��/'	�)����{k�8ʶ�^,Z�8{���N���V�]�x��:����_w�a&$;�)�	��k龩�����>ߘ#_�� ��I�X{z�;���������ۗp;
zN�]���%�偉��~�ٻ3�3�Ƞm�w	�s<M{�zU�oI�U]81\�t�R�)���� ����NZ���W��\	t��yn3+q�� ����z�|}��CX@��d[�8~o^�&(�˅3�n���TH��<I�GW���,���|�#���lKN+.�Mk���vLY��M�Nf�1��01�����J�AX�y����	�����"��t^Q׈JO����f�@�^�e�[��D�c����$�&55o�!��Ѯ�/P���盋?�����5�ɱ�|�E�:�=�_��ra��Z9�t~G���5c���K-�,h�eDHk\r�����-�&�i:m���!8��^;�K�Gu�b:]�t�@�X��a]��y�6W&� �ͽ�,z�+>���]pdƏ��6�e�3��:,�S3`��s����ƛ�����[7�SG49�N&�º�(���M{O}��5�����ȟ�ʺa{�t��)W���v��K�-+P��������M�e�h�xz<j�΂����r�'�L��U�c˝s9 ��l�m��q���ݐ�imQ�a���� �b�($���t��.UI�s��Y{������{Y CN`�O����BQ<C�����T����F���8ɨ-���&c����BƸR�,
Ql]9�@���R;� �Y����K��s��n?8U&_ x89L�8�	V���S6p��0ͧC��mf�aoX�@L9Y�Nm�V���U,:�2��2��r�U&Io�%��<9ˆ���A�⡥D�k�h�-HOL��6���q%G�Ewi��n�'��잉K��?�w��P��\�����9S~F�2���l�[�M��0y��y�5?�G�2ot��C���hdS�c$o��DPw��\��4�f�/o��H��n�r�m76���>r,z����.&1��������f$����#2��=7��꩓�����<�*VX���Fz�n��bz��^n)����8q�ຫ�ag ��*o�HE��jL���x��m"�<�`]%ӾYP�����2}T_���;jt�N>Aϥ/��V�v4� �W�J�B�x�6�QrbH�85���%ͬ:������N�,iC�+8=�@�ᷔ-������@�dJ\�G ������Ř�!v��j��\�:v��1����9][�����D��������z�v�u���"Tkr�I���+��!����݂�+}�7��r��70����ڗ�ɠ�XC4V�5����k+���Pp\8�V�s+�i�G��_8�