----------------------------------------------------------------------------------
-- Company: BINP
-- Engineer: Epshteyn Leonid
-- 
-- Create Date:    09:45:30 04/19/2018 
-- Design Name: 
-- Module Name:    FindMaxAmp - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: v.1.0
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

library work;
use work.parameters.all;

entity FindMaxAmp is
    Port ( In_Data 			: in  STD_LOGIC_VECTOR (127 downto 0);
           RegInit 			: in 	STD_LOGIC;
           MaxAmp 			: out	STD_LOGIC_VECTOR (9 downto 0);
           MaxCellNumbere 	: out STD_LOGIC_VECTOR (7 downto 0);
           ThrNum1 			: out STD_LOGIC_VECTOR (3 downto 0);
           ThrNum2 			: out STD_LOGIC_VECTOR (3 downto 0);
           ThrNum3 			: out  STD_LOGIC_VECTOR (3 downto 0);
           FastTrig 			: out  STD_LOGIC;
           Trig 				: out  STD_LOGIC;
           SaveTrigData 	: out  STD_LOGIC;
           
			  Clock 				: in  STD_LOGIC;
           Clock160 			: in  STD_LOGIC;
			  
           Reset 				: in  STD_LOGIC;
           ResetAll 			: out  STD_LOGIC;
           Error 				: out  STD_LOGIC;
			  
           test 				: out  STD_LOGIC_VECTOR (15 downto 0));
end FindMaxAmp;

architecture Behavioral of FindMaxAmp is

begin


end Behavioral;

