XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���6Ee�1#P.a}n��vڽ�e,�5N^t��1A?�[=�P��c�ɳ��,`slP�_k`#��z1tu�����7�4➼waA\��q���O�P&���%ܽzfd[D�k��n�Z����a�l�#-����A�z)F�귵��LY��Y$�G.),�x���k��6�M�ac-+XYPRInV�Ғ6��7�e_j��E�-����.�#�H��|W���Tl-=����W�x/.��VSâ���	��]�� ���PK��~۱�n�������/1�T�=��hѪ@�2�N��pF�:�h$z��E������@�>�7F�R"�����]&Y���/�Re�����6ykB����u�\�߷��f_ȳ��c^�~1�-�X�@D?�iq��8[i%y�Wڷ�^��e4�RN��R��\b����|����i���L�R*8d��mLlsԞR�z�񭷆��2xt҆����Ø�}��>㑫��eB���	1%P, ab��A5	H�J5\�b��Q�ZI�SW��,��e�#�4�Pt2D�%?Yy]�S�[��¯���J[��ՈK�{)�1�Wq��V��,��uٟh�[5��PG�Y�Ý`���~�P�i3����-tK��/��%2O��m�K��h�O��k�S�v��~��e�@K�	�19��M�A�#_{%^7� >M3
@����$ެ�"8��r��N奉�wx v�J�|��򵓶�[�(��J�Q��o����6JjC�^_�~	�Ϝ��XlxVHYEB    1231     7c0	�v���^�����tz��D��l8Cß��8�h@�>qV���d����-V��L>���Am�� )(.�?'̠���H���6�|c*>�1e�>FM��vZ~���Fb��Fx�O���G^Q�>�������Ur��]�V�L!v��E7˛�cֳ���~��c ��n)��&�w��C#-<���j��pC��xS�-,�t_�x+�y�������p�6l�++٩P��	6��}FĞ�y��I}n���&aFy�@�R� #	���@Z��F5���ffK�'u�od ����e�k���O���]c���7|x��	�R]����'�[�r���"����M�(�h�H`��*���V���K�瓜/U���P�0�)�:�C,A�dS��@�q獶O�?�ǆT����D0�R���@L�ei�Ԓr�/]��$�̼�� �+��GOZ�������˷��T��dY���7M����F%"�tdL�8r�WĴ�M�yJy��xR(�
���Tp,�|(ఞ���>A�6Q���R6Q�n�Ug������B��k��*�ph~��`�r~ǠV�s��*UL�G+G@~	��%��\g�z��7Zg�n���v*�Mr7�����`���jɒ�������+Q�c����)�&c7eO,�� #�|�����#f�M5�3/9����a�V5	�9{���W#������k�bvغ-c�w�+[wϮ��|R��i��9�܏�j0/ѴB��]飳�J�ǲ�Ty�2���"�-T{B�����Э�(.\Y�����y�-z̋�H�#��27#4��7P�Bv(�X���OSMu��KL�ϐ0La���l��*�Eqނ'���#P��@	�2�ж�Ufl%,�O$�ƀ���L�:v��6�&�o���va�/�K &A�y��Te,�cB�����(��7���
Q=QO�4��t�����:������2���JL\@�K����
��Z{�����Y�����A3�;`�%
J�P��[t�5�V]��Ƿ�n�8�oR��Qp^ܵ+����xV����o$�ڿ1�Gm�.Eь���s"m� Ri� ᒼ�a�Α�K�*�i�~�����r�r�C�**u�����~M�.�gt�?S0e�%��o!k~�ȍ��������-�?	�%��K 9��)OƉ�Y�l֚3W������Q[u�Gԉ�����H��)���T�le���V�*pl\h1��yl�>l�7m5O�T�=����#��)�Y~h3<�X�q�$0duK�H���#&�Z���n��Z����uL)P:kG�q��BI��YG�wt���� �'y)�Ef�PGA����>��hT��c�\�B��w��5�_פ��o�V�,zݚ�N&l��z`��F�r��P�Fk�Ɠ���{e��͸�n�hÀ��41�(Q��"�a�瀠�w:��?JQ-� Z�
F*<�������9�n������Tɞ����q�ܜr�A���\��<�6F��L.k���K����V�
�ԇA�46��7Ꭓ��.��+�޿��+J@�]�e8��&�@�`[5��T�`�����8�nYgR�a���������#7�x1��~Ί�0tp����Z�3�}@����I���8=j��ꝼS�z�����x�=L�8(�w7!�}�e=,% ��y,��%(s4\���w��K���,�����aB���y�8���Y��(^�5iP��'�0��)�����Vd�s��3L��"m�w/^�z���K%�^�\��	@�����C�?�1N���!������+¸��}')Hb���E{0��`��o����B~��L.�n@�h�u�|D6���8��1����4�o��7����߄��e���6D�&]0ú�S��)U�����m�H��_(di-wO�ozPt��qЀ/��,������"�ꋛ�`D���,