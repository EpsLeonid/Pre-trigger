XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G�&�&������X�"|�Zm�<��,i�alRs�uX�N`�4/�Nw��$�Z�8�@�q�2�|���
�n�B�*����E	����T�Xg�z�g��� ~��r��>Q[aSE�<�^ӫ���8]l�$��$���S%�����8�˴6�O�ؠ�#X��V�Wb�����˛���b���pG�m��k�g�͹��:�A�0��B�������^a>� =�n�AR�Կ�T��~l]Ǯ"�f<�|��y:�}���*e��u�{Y뜘�]zQ�ï�c!�+������a����Y��#����yfM�͛�T�ރ¸�M
H�X�V�A���շ�c�!Ogr[j�K
�9��*C���M�	][s1�)��]�a�&��ћ�=���Q��7�iv�>J�d]����d�v���M�R=�#�d)'*o���;q�q4�Kh�fː�ʐW��if����r��<�����m)�����)�!�}�����D�
a񰫌����m���7�g\�=��Ai�I?�pM
���튠�+��+I�� f��ZK�pE$EVY���E�4�"]��³�{1e��v��]g�8��)� �L(�3_z������Z%�8��$��ꜗ),�Ќ]�Eo����T,�ɶN��A�[m|Wl�w�;u���d�lw�{��}r�$�w3����>?��[�fP�c���3WAU�P��H&�}��Aݝ�o�"��������A��rA8���,XlxVHYEB    47d6    1030 �=��"8& �`i_��}��J���R�,Ǿa ���>��y�����Bv���x�r��v��E4F(B��#��p�s�X��o���A�Z�>=��v���G%���|�퇏�v2��L��(������q�}�,w�V?�@?$z�%5M������ֺ���1"�xE��)��1>�	�W¦YPlVN7���{EB�p(m%��w���Z��h��O�M K���"�{B�e��6�T�z�N7]NH�;���O �a�u�M\d�/u�"!���96 CpǞ�L-J�tD%�q�.\���[��<|�3��b�UT�3?����5�.���	�"R���A��������{�v�g}�:�9'�iu��e��`�9���~s�g!BP�u��Lnn��
#Z�o9-�6��_�q��P�<�fD���"(�H�Ĺh���3�4yJ�)�ū5�Ò�=��7�w@mk��&�W��v�8�ڡM>�eyŦ^���C��f0��f�q�W����O�l�ԒR���S�o�	�����zA��iM�����YA�J�P�1/�AZ�7X��cb%�*m�Dw�q.1O�T�x��94�^^=7Z^��A>��C��R*[����ղ)���c�aɩ+�y(=����O��r�y�(��3�~(4*,00���@�h�{�l�s��1ƮM��#��Kzu�'���w����y�����q���.p�{����׵7�q�}��T�i���z�N��"�%�)׳��� ����pc����
^���^���#�ȉ�ඥ>�t��]�8c�A�pP������b~��4��t7kH����II��G�ء̋&T[e��y�EM�ᨱ��Y>��E�9��L� ���Zۇ���Xs��h|LY�2��Y���r��ĝP�7�b��҇��ċ��]_�_C '��˂L�aIu>�T�>���x�}Jv�^(�0M�����m.a
&���;�:�I��/�:�A�
z>�Izj��i��ۉ��u6狑J�ӥ@�3OZ��]X�	G ��.������0��`g�̭�-L�~`�G�x���N]?�;�ɶ��Z�2��z��z!aSr���#�v&;]��A,h���"g�	`��3ƻȟ��C�
]Hs&`1W��{ޞ!c�\4�ظ8��x5I{�{�=lP�-w�l�[��x��T`�ϲ�3x�n �O���`r0k�:c.���j�N��$n7v�9�=�
L�&��t��J2e����2��\ ;)��Etl{5�'�}�Y��ز/����>V4s���}ݰ�g���P��J�'����Z �
4ʎ�l�k���1����c�E~2SH���}ϫqP���$�=������J���ͯ���
�	g3&�W��-A]�a��,mg���%�W">�C蘔ɮ�B��y�U�Up˳jy��j�<��=��qx�2��R�AFy�U��zc�wY�C�c���n�R,
�W��Aoq�O��x�ڿ�Tp[�A�S�[{����ՄS��6
w
��z�r�@��z4����x-��\;�u����Vp�g��"�}��k�}��c1C�?������)��c/H:�S5�7�}��S��i�@�	"N�}�����)�(
%kP�p B9'�����y������]枪\F�t�i��o 7]a@��f�*NV������+d\������i�5�T2$�2�N���$�Ck�\�h�Lr~�@��a�Pay�@��������)j��,	sKu��Z�StҴ���Y�wkF��T�o����f�"ic9u��;]>ک�{�J�f8��e��] tE{���v�Je��T��L�hi;F�#L��� %���'�蚜��Kf�V�UC��G�g��~��V���1DϚ�e��hNRt�Gg� ��Ub��t��,�?g�3L�q%�6rB�Bqʟ˔b����;�Ab�Sd��Qx��v5B0��:�5����'֊`�l��!'�;���^�1��F�Ɖ��mհB��b��T��!��K�*��-T:�*�5&>S� A��؇6�(:�J���.l���׹��!z΢P̾v�
�̯��D�����Kr[��lj(@_� t?���A]�G��u�!�7��ThI�f�+*���(�l�]������g6�d${��}Ui���6ԴA��|u(cۄ�� 4D���b��Z��x�╎�,0.���*�?�)Z����ko��H͜�.�LĬ2?��iȻ��(3Vظ��%ʶv!��`��2��x9j�;,#��۬���~���l*�Ρ�y`0�S�B
��J3K ���7�ocD����Y�)�"�Vf_
��k'ꠉ�St�"��J$w�S4LG�g����,i�Mv��*�֢��oD��FYlAFĳ���E',��wO�a�Zš��q���$т╪ɩ�'u��7b��*�n��L]T�'�a��}5E�y�x��k���_�P�v�#�+���=%�X38G� 5�Y��K0j����"�Q���߈h�u��$5���q'|wz>2��P���a�@O�p����G�L���*���9��9��M�Fh4z�t?|�dm!�gg9D�H�Fu��i��c���r4�=�l��HE����vdZ��<c�/��bl]�����?����W�ƀd��Vr{�*�Ԅ��=p���&��D�L����^?�C��6�y��<~�B�=�ǀ���G'�$�65#!�k$�`k�}�g�ѥ?1�|x��c��<v�$������@I�v����K�����`��/na��-_�Q3���̌��->�T@���Vv��Ag���L��W��*xܔ-=�ξ�8$p~�-�q��F0[�`�a��Sd��]���������� ��� ���,�2�x���y|���� � �O�D�b2��Ѭ�P}e�����`9j�и!'��H[v�V��BaCҗv�:MU3?�$���C��kgrYG��_���}��흂�p/q!2s��a:���q�{|`�x��}��"�U�3��Ѫ<�p�K�Ɖ��H���T�\�L�LȮA�/U�1	��)��E�)��g#�c�l[�eU�~��#�QcΨ�0���<�����ʈ���\���ɸ�hȬ�0UYR���5��_�3��S��k��P4!�¬�&U���P����ή�>�u
��e-�U��$��ټ৭�/�|����n&I�����ڏkZ}��~�)/����\��b^��׼v�i�J����5�cY�a����3'��UZ�H�ԭ��]�����u�ߕB.<�5����x��X$O*/��x��qxGެ"V;9�\X.DJs��f�i%��7��!)< �.����x�-4ek���E��xHz�
��'�*��U2`���s���k�[�4�[�H�s9-:�-�a�4����-�?k��_阡ϒ)5�y=�3,�����8�����n֓��C��@��x~,����v��)�N�̠cf�30� �@�;������A.P7|_B^�e�ϔ����Y��q�IM��b�D�IZ�Џ��Cs�����FRk�__������II��#=������Zb<]P������z��� �JW S>�ز��X'�F�P�����E���}"�	V�,�������D�8b�U��#pp�_�V��&Y�H���c�*��Ba-��V��Ie-�]�ƞ� ��'���w����T��MX��k�;`�����e��	�B��m�#T$����X�)���]LT�O�H&����T&��A�Fu�7A�h���'ߪ3�K~["B�� ��3�O�$��_��²�-���]��'2���949�Ȧ+�[�)]W�h�!�3�q˧���|Ѵ)i����P��"���2�x/Ĳ��c�8Ϋ@�)���>�x�����ȋ �/��Ⱦ���ɏi36�	����:T(��\]�?l����'��=����$e��~t	K�ϑ��Ș��Xe�x�<g X�OUn|ˬ V!*��Qd���{��`���X��:S���W�H#&�7UvP#�m�e+9����-%��D6Z��Ǫ!�K?���1�rr�����ny�