XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;H��^��J)з���*��g\�������;W�F>�.%��]e"\?���!g2}(%W]TA�e��2�n�.�ԩ��F�y�.�n	7����6S��:�>DCG��~����d�Sw��Z�����m(�ޱ͐%5Ĵ�WF>�C����P�3���=G�K�\"T��^|L,	�wK�a��imĄ�)0��O��Y��ٱ`#� q�Db}Y�x���O���9�ӣ��Hb�k���Nȉ��/�èB#�=���Z�5!VZ�I�\��Q�H�,g��=j&�J�����L��G��|��TA�[ƶۤXyڴ �0*C����$-�UO�Iƣ�J3�$|����)�跷���ޏ*����8Ϫ���&�W��_�4S�e��5���C��U�+�
��_]�����z㝰5�)�	�⺍���,%��=R���M���S���L ,�T�l�ĻiW �|�s-K�_�h���yĈ�d�����Gߥ	������R2ʖ�i�H�s���r
�L��+$�����w�Ќ\��Iվ+�Y�A�y�u�t�E�}�޺�����J����P�,���7�"5'�;�CH�ݖE��>������׸	Ue"�P�2i�.H����~$[� o�K;������]��n�&�S�.�I� 8j�.)�!�,�L"+-t|��z���si�aN���%{8ih�����9�]\�j���~���1�̬���vD�o�x���L���4 ك&�O)�XlxVHYEB    1854     8a0��x�1bL?�z�nƖ��7��Ȟ�'
;y�� Z,�`��1�>'�~;�� Dm��we�p�K�U�	���XOy̍�vVl;�_#~�kͺ������c+��mQ���z=Q.8q_h�;�_��9)q���&���o[x6�p/�X��m��B�|.��?<l4�do~"�3X��ǜ� �g�Q_�^���ٖ�~/��C��]7��>1�گB�`��׃�<�!w2��"7�g��[H^����K��̯��q/�葬��ȑ�5Q��?Hy�3vp�Q�:�w�uhTH'WT����&�B�JjG�� 8T����Jy������5�.0oң�*��~J��'<�M�� �M��N�Y���c˿�_�@_!��<bO��Eb���V�l���Du�?�/Ǐ�RCdU��<P�g��:�`���ͻ�H�l�{5�k�#��w�J+J���M�r���! �n���i�V��/f\�ot��c�9�l ��fnpv1%25`֦L�dQn�� ؞>-����h�`�(b�s�����,K��OW>rr���N-v?��)���� @�l.�L�'�O"����C(��
��,��w���>��dwN;�~�)�(���;�Ĵ���|�5SΊC�������80Y���	;�}�� ����,_^��:�R�UŦNȴ�p{���ATĐ�W��L���O&:�C��e(�-t��!bw��˂�gd�ž���:V��tn�a&JE[d�h��l�P5mٳi��(�{���`���B
{��m���Uw��L�U�Sc%��WTU$�쾏R���cEL�{>~U^���-@'�tJ���!�����w|G!�6>��,��7U�|�cӉ^n�i�q9�蜊Q��`���Y�����B�w�8O����#�g�7�b�9�}k���!i9�v�`TN�`�8�~���y/{�2����!�QWb��k��˴��=�PF�#�NS�)s���s],:,Tu��2�Ч�
�ڏh-#rl���I���*��l-����b�{��^wx>�!�C��4^t��52H�U���Hx��.%�&���q��{Ɣ�Jq|��b���]�֡�d;���ȒnR��J�I9E�x�8[&y
!\kt#d>�̸lRi[�u��&u��nY�T����FЉ�f�0�r/�F�����d3D�������y^��ׇI�H��E�.���W���\�	.J֞N�wfs-���޻�%��W�h"�}���WƷ������P�{��H���Y�>���}��W+� c�G��HO@Q7`6|Y�^�Z�ǘ��eyv�ɀ�����Z�����d��1��eFRGNG�>r�VF��r��~��c$�&��2��/{�QCkv7��]3}!�}�Wh�
�9@�CC��`'�$���G���Hm'�R��K�A��+A��LU�RNC~fSpl�
�(������mԳW� y�8*�����^�{f��)0R}��@Q�{����(ׂqa��}�D�dO�-�|�O:��PW���j���$U���+������E�����c+�Xyd�iCD�?4��S;nƅ�v��W�T%���>NN�d�Z\���`Q����T�th�bb!����HLX�����30~��Y�;ӎ!jb���.�c'E�0���"����T܊"����
�2|"�|K`�Nj<��kD�8h��fPD:GxqSE�o��2��`&di�C�!��y�oQ�n�y�י���TЛ�Cf����Β.�[�:��_je�ڄ�J��t��.C�����ge�b��@sOVƜ�{��G�*����n����6���׶��kj�/�I��0g�,�&�q*e�����.� h/ |�v�i>¦�����/��zJig�P���T;�+�O����I�99�;f�I��mX{fMX�۞v�~2{�(�\*�R�ڐ��,ȖP��.��R�L�E�Um�{VIf=^�Y����<)��'M\M�@������䓯��)B`X�����������C�	�?NU�(]�=�c#"�&��˧��#�wWǢ���?76�a+���u�\1�ߒ�|�ѯ<�\|�o7ٖ����2�?�"�܌3d^�Xs�Dt�'k��io���6�K��~��'1(�������)�ܹ�Œ����B�q� 1���%�0�ruB