XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-LcI؆+�G�}0�ߠ�v[0Av���%�XΦ��5{�"����,f�ކ�H�ߚ��C��tu=�E���Ȼ�7Z���L[E��I(o3���d����/a����d�`r���@�ڜ����~:��xwq^kH���~��Ǯ��߿�1�;��?I^��B��2���g��#��Ǭ��?�G�cj��z�J'����L��x�x_��w#�n5+�f�`�䄁��]G/�+ԋ�_"p�n
����`L�����d?�͊��kky����*�&
0���Q����1W�ͽ�_M�DJ�L�la��JB�;��&��/����c`��rtC���`C{n�y����%��ں'��(	f����1�ݞ �'�FL�:a�s������9YQ�"y�Ct���\Z,m,�͂��������b�HP7�;��=\�+In_9=6��: r������v�0B�^�4����}k����k�|i���鷶.Ss�'�;�F� .����h����z#��F��>�g���{�@C�J1��Q梩l)3JG����Z�3��."�i�}JDъ�ֲqJf5Q�D]���j�T��'(�"�%�ݙ�A���r��[�XU���)��B�����,]�'B��@x��,{ϷzU I��}�p<�~تղCe_�yW�����N��QC�%|W���.7 �U�Vr��3d�6�W�^^@�raܞS-	N3K!uq좰���pQ#N���l�XlxVHYEB    3f19     db0z�I�ޱ�Z��0+��&[g�l]YX���4H�GTSh�k�b�]��3\^|�"W�ga�DUK�|~?_
.��B�{l��J^��������Z����t{2�ģ �2	��rc�N]ؚ?��vU )�L��ad=?�P�mz��b�t�k��Y2.JkU�a��o�=�0 �~,�s� �P#{ˡ�8�ءk�/DU��F�r��=m��ei�7ژ9#d�`K}�~[��8:��ж����	�衠0�jQ���D�|��|�Ǳz�]bt�',D�÷t:L����ܴw7�H����u� x�s	�@����WDx}�C����@c���m���~�V��o���ɽ�0�ŠX�{�	����-����(�FԱL��Z����~�E�?�g�/T8��������i���#��vbe�ɇ$�\��k4sm����V6�WjK�	T^����j	���5 O�K�ذ!	x��Q��}4_��v�7�����ߩ��phg&��k���M��巤��~�+{Ǘlf	�kS��Fe��־}����&!�V �>�l����M��m��#�8�n&V2*��03voVx��N.�7��igh�t7�(�ʺ��w�?�!`h���C4�[�'����R� r�0�O�5�;�a�e�����h7K�K����xm�C�����Io�T�O�jK�*T�X�wD_m6h�~7�Ж�+j銛�����9ûx�_@Q[nLn�kv�s2F\�����ß0h^��W��de�+d�����G��=�>�"�X�9�B%Av���sX$	%�f�s����<8e?W�V��	e���;1ؘ{z�<4=�ǾK �gn\_��[�K��[O~:P�"����Cu�TVB��
��.I�o>�@����� \�ސ�gF��O�m�LV�,�o�����g��]�Vya��N��%����,���gz�B���f�\
�4+�d^ ���ц�3M�Q-�f�V;��s5���a���g ���u�'Ͼ�oF3�Xx=��;�-@�<�<����a�j)���˶�떸��"(��eML�C�c0�@%`^�/T,Y�1"P��~1�`�a�ﱅ�?�{%�E�*w�I;a�.�Z��y�t*���V^���+���+�G<�����ŕ��v��Lb�E��a��j� /<Z�rk�U,EJIع5,�r,�S��@[�谦���Z{߉V���Ǌ@ ���s���J�z�����$L�'`n[�# �l[���o�x�*2���\5k�[ ���������[y�
]2.
�:�h���:� �rpt��\ѣ��Y ,4%Q�fVui��X�ǫb#6-Ŋ��\�3gF��5�$�w.�J_��M�~��
��J-?԰��x����>�w�3���&&2�Mv5D����u��06�ƶ9�
Y��4���0����2.��!y�B%�:�s��p��%.�H��WN�r�*� *��Y���nƊ����^$��jN��_ �v�^�J��Qܚ�Àp|o����X�g�]A�4��s�����w��+@�𗱀�J1,迼تX�ﲵ�N����tV�:R-�L:[9`��_b&��dk͎�~ɐ��6ُ�(��|�ˁ�g"WQ�)��ۨNȾ��9gr��<c���]�I>��$0�'������/v �B�T�,�����0��+px3��L�c��N���)���7��H�h�T-��<Py�˚�I�A�����<}�ð�S�P������q�74����{�3�is��Z�}�朦���5��b�#̷˅%�hh��q�o+�iT�tOY�)�+ݠ����McՇ�#-.�Sۂ�L�d΅���5s���W/���Q������$�FaE|K�.��ffa$��	�9���K!FYp� #Ϟ��U� :��=٘bG��7P�hB�±�1��H��1��e�S���W���o&�PQ_��'�o�k�E��+����1)m�(NPZ��M/iG]HFN<�o�����Rn�ûtW:��C���EP��$�&���)�EA���rb�9;�<Wo�jO׆���pw�5��#p�gL}�p��_�(msL�=BO�w_�qiF��*p�	���=Z�N��Xv_fVe�:�#��Rv,�� `_�hG�c%�QC��� 0}�����1ۀ<����Yb�<��#���<���iƢ)6�c������v �7��V��hj+�i˕��j���yZ �)
ʎC�A��T)]�2`�Zs1�\0�)�3LW���)�4�	�CP#l߿u]o���F��r���G_(��Hl�Uc�)�ڣP��3���f<����4�r�&Q��,��ÏKB|)Q��s��:�O>��[���T�ތꁿչ��ʌ���M~�2�$��M��YeOA9�V^�� �_�`>�gǏ���G7O��z����tA:��ed��$��~������+V��`b�4�ѧ�[�K<�,���Gx?��l'L����<��I+؃h>�I�)=�D=�0%����m�n��Kk8!�W>���'���������6��ϣb��Ɍ��c"W�o�d �AR3��iK�=��i�[�ݚ�ڠ����r@*D�9�&bƾ�p~�D`i�I�9N#\����[��1��$A��"N�2ȍ��e/p�Xibw�}j1�+�X�$	�����ch ��%���[ԁif&r�&�l�Лl8��K+�1֫)�i�$)ٛ�ٟާON��~o�4�v�e����1!K�Ey2,��U�8�|WOp1� m�A��S�v��>�w8v}[��ٶ�V��;\b�1�T4�J����R��.�:���N�m��^j]����4��[ �{�6( $�W9�ٖ�o�4�B6R�Dqa_����D(�-�"�z�:Df���h�M����xԏc^j)8%�[�:�!T���i>��x�� �!��a ; �K[���>�7��z���8��R�������Ԅ�P�L0$��EK������X��{S� �د8��+y��
��#aN_�DU�n```��M-���7���F_��r�q����%�X�n�U-��plik�A����� Ӈ������E��s�,ϩzc��Y�k��?IOP�Z�
5���l����4&�^q��(a��K�
>��۾�i�6�)�8k?+_ҦBy��A;�K-�(q�� �sl
�YU)$�^�V�V �~�%�?UH��=��_9��yh��cc���Uz�rXCN�+L��qD"�@W�=������c���;'�/�9���x�Js��$��S;��$����en��d+��(��Y�������%�-��.f�%v�� �C�k狗�i��d��v�G>�:ğ$�&:iAX���X(*Xې+2�d|C[pA->6:ʮ����}5�8�Rޛ��~�QN=�WA=)��FH+ET�5/#�C=͵���U�8o	Z�@#�k��|������k��V0��