XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���]��R3g��}�C݉����Gi�����E��LE/����H�J%�_�=6�b@]��2屒��r���6�&�
T�z�Ä�{@z�\%� t�*����Ni��vjh�h�5w��}Uz��bO�`N^J�ס1ww���i@0.�U?-�»ā<��;��y+�nVc5�;�sq
p����@���0?z�����ð!"�D�+��F��>���A�p?F��e�-	���}4\�7+ԍZ�=�B {ڒ=e�������� W��H������!$�fz��Z��vL�V���߷کk�׳
�ڝXLS��$<�o�ڪP�$Xp��_��
c{6Z�J�i~,��߾D�_>�--��NX���*E,`T}������0|��L{��ۃ(����ųx6t�l��������_����l�_�U4�%}|�2Y���<����U�!K� ��3����jIDuC�NeZ4a�ᓚ(�W@��V%�i��Z���7 n9e1^8�SV~z��#۲���F��"����^�S�����
�I�0�sH�<V����0�)�Y�ěRѨC�h���C�� �9#�o�]��;O0f+vP�z#��l�2N j�&��Og�O^�� E���[Q�M����]7>H��=-#XD5S���S�]~� �H}����P�})~T��}��}<T�#����]�<M*I�BK���ŉ�5�&�GǘS
 s-�?G���_4
��j8�7�_(��?�ϽXlxVHYEB    3f19     db0�r��2
6�D�
���}�c���9�� ��K��3��&
�nFs0yu���̶~���O;NMvֽ7ٛ!��d15���n�`���K�*!��L�wZ���MvG~ٱ�g��C��1e�D���4$|{�99+�9�E4�S��Fh@�
�������z�m������|�!Aa��0����k�U�Ч����5��@�+H��������XQ�0r\uO� U2�+g��H�@�U#�֘!��:�Y��\�}�:S�Le~8A[ڐ�Kx�l���C�r��'C¦���J`P��T�X׹S":�Y��f�h �DӖ��4�b��/v>jfm�����|5vx �PW���oFa�M��kyS�a}َ0H�0�NL�_:�u��z��I��5h�G3t�y$�t�R�$~�����qd6�v������W�cYǡ���t1��7Gn�_Խ�ja6>�|;�~��@}����gj�^���wbb�%0O�ZٲXМ��Lo硐�-8�[�u8;�ޢ�1��z+MD�S	��R\�K�.k�4ֳ���L���se�ǝ2(	�	Fc߱�Qr���V�<H����µ[P���?pk(5�6���$�zO
GN�&�W?�y{�!�vyO�Mb�U���.� {�)b-M��+�E��/�TkC����6�?�dtuζ��p��%L�ԠV���ۛe+��_�ج�#	��LІ�)��+��5���?�y�BY�>�0wS0�g��+��j��|t�cM/� (8QZ�ȓn�痲��bXU��r�v��� �5q�En����_t�a�o-��D�Lz���x?G��!nv�?6�iA�Wave;Dm�w�I����5� `�eG9�|z��c��6����!2
��ef7,c�����@ueG�b�>���~��HT�a�Y��7�۠Δ����G�{#E�[t%���u��gݟ˒�m[�y-V�O� �g�3�{3�.����ێ฀VD!���/�מ;ڠ������1�]��E��W2qd��FA���I�P�K�Q����U3���IT�74Q�+��]�s=g�3����/�L'��i+�Q�n�Bi(=�)y�5Gӥ�3�D�#.:N��^��ѧ��0T���B|X��Y�����^E)0�>0_+䍳�d��}0z֕�_�cX\�~5�(�8�(W҃�Pg��"���B��J0���'��ScT䋅�+H��3����Y�~D3���K�o��L��=�#K�L>z�V'�>70!�.�vʠ�� C�XH�q���(����ہ���ˉЋi�uu��O�3��v�Z�,Y}B{s���;۲��v?��Z��9��T�*��6D:�=H��m�,�੉p�U�]R�҅�Wξ��9l +��(گa<*�ڤ#X�� �Uw�:[��]�ɕ3�ѹ@�r׀��h����A�俍���_?Qf�h��mL��ѶC�lB�{K2�j�q,���Hi���V�c#����u'��ͼ�2D�@v�<q�V�èG��#VGi�q	+^�h�]�~�o�%oxR�ݳ�)4�۲�IӺ͎b:B����7����������>D��-*M�����@�����us��3A�p���8�`�����%�M��?���I
��x-���h��%���#�l���9���w3� �5��a��Z���rD�7���n��1	wc��oS�~!@�(3�.� ���gr�T6��ےU]ǌ��?�"���:��g�{h���F��T�yE'@���
�kر��FYҢ�呿����u��^��e�����&��E�a�Y�TF����*/��k�g\�y�\W��O r�$7|�Y�����c��-T_^��w�]#͜jT��d	;���.j{:��P�{*}���g��d2E��QG�c⼲�+"'e�r���8���|�p�ޟ����B���tTޫ$�Sb`����YA,�ή����"IQvH��uk��>�0=(Լ(n��9p/�n�<�@��"��-#a,i�*��Z����쎾��97f����"�i͇��A�;2����Q,�L1� /����7J��pf�)��l2C�Ϯ>{N��k�����M�P�']"J9��
��-FG�;�(+��[���.���}?���
<��M*0��u�á�W���\6�T�v�D�ߔa��?+,����DݟF�J���c�"�����0@)"�O�iIdSƜ�����I��ۛ\��Yb���=0#�J�,V�I���dyn�D��R��1�_S����DM@.#r�͜a��֐�����"x�4������sdy��J�i�F���yE���(��,|��)��y�WY�i	T�[���]k��-��yx
x����/<ʩR�h�`�K)����u�G[��ۥ�*�x���D����~�KQ�եߵ0��3L@�P�m���`Ȅ��G��n�u�S�����L�u�?7vYF���_ ������5�2/���&h'K+ˤ�������8�!��f_��U����'(������f'h�����,����?����d�-
�?�H_vi�/jH>�6���5�n�}��hj�d�pa������ެS+��Q`��}� �z����r�T����/3'��:U��?�A���ģI�u9� !EM:ƘQ�u����������~�T浘����TvЛ���Y�̦�Zo.ع����;;,_5Z��ḅ~��g���(퓘�.��F#��4�&���&#,�4�}���(�k�uT��Cd�V)�_憧"��Ce�dH�D�*���}]o�:! /���5�mI*���^R���Q9}�d+�~löf^��@`B�U9e��!~A+��N��D� V�c�d	z����r+9\�s���F��_���'dl��:cj&�^��h�C!�̭��.�^�K1+5�[d1��P8J��� ���d��a�I�*7� �Z�ȌR�vZr��ip�j�<sUB��C�,��.��+��ys���Cq��3׹tl�\C�ʂ�mr-J|��mV���*�u-l��H
�����tԑi̧"/�g�&��c�=O����S���[�^���^�����]��q]�"d��h����#�b"y�;�Ӟ�͎����1,��#���n����#�+���i�>S��9:��\�����L;����u�8����C��>�v�$�Jb�C��p�_Y������m �=�ڲ�ne��_�)�`��i�^�]��beMe6�]�O˂�z�PBA`���G���G���iqX'3�#P�7|�����n�3 �)���.��/*���V�/�9:�
Ἰä�R͝��c+Z�!>�%4��֔��'��/��$Y_ۍ�?{~D"���1mS�Ɨ`X5+��Q!0��XEs����׶ZUcW=�'2uI��b��e�zގ۾���(ܗE�iV|�4�