XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���%�։0��#3ʺ��*�?��ȉ��t=&;#�6�-��K����*U-oZ�dA;ZLN`LA|zRH�3R�5���E�ZԄ�tD�#Q����z;El��Qk3q�c�������n���7���x���KB�[Ȫ��(z{`�.k����:�AN���]3�O���4|д��(;��l�,9�N[��p4(��XBbb6�T%Q�@���k��#�E���ƽށq�ڀ.��@�GoĚ(Ћ��9��ǺH���?�<a&~;d�o_�REI��(�?���)�7������$/*A�Y�a�y���4�Zﳟ�=~?TZa5���F7b�\�Ci���'��`8�� ÷�8@»��^،�GC�9���
�
_��w��]��6Z�"�ڐ��Q��X2�;��/c�m��PA�髝j
KɧճĚ?e���闫�^�<(0<�.RG �����e��㣠�K��<e����V��VPy$�ޝ�כ`�RxC��L�$0/g�L��۬�Q�)ϙ�:*�r
�D��aY�S�P_~�gė|�ųW�|�ɓ@�\�\�9V)3 ;�)�3��<k��I�X��'��	�#V8�U��=?��}�j��]�b�밳��]�����
��C�w�S���̐X�h`�4ж�J�}ϟ������?�.��?C�h�CX=�3(�ڄ͸Ó��3nN$���ݾ�>It�����X>�>9ؔ�Ya/o4����<���7�%�ͺa�D�w{.�@hӫhmW8�/d�XlxVHYEB    5f5a    1490Fj�Fl�UP�lu�Ҽ����IW
��V�����/)�w?��畴|���	#��5U�2)/�<�R.�ϯ�y�N��p;q�K�H��/��,Ga���A�z�[�=PIuFv}!�}��q�%�t�]�0��7��K�X�:F�ݝH����_ԛ���se��G\��]Wzm�h��U^o��}9ǁ*�J�4p�'�#��=�0�o�3:��|N<�tE1�1�����	��O0�$=w�kr�Ф:�\�ɱ����u��F�}3�I�L[��Y��;6�&:
f��[Ny1�>M?��m^����ց�O?���&#;@	�&�%���"u�^�g,��/+�%��ou"��G��9v9�[0��%Q�[�ɋq��Ӏ$~�Q[i�kM�H Y
��h�v�9�y���劝BJ֧�.��I�4sￛtG����#n��������:UŸ�]�(�F���(3���| ���%j���7yc�oﻚ
hќ�{X½l�=���&�}싦(���`S+dY��qn~\{y����h|gj[̑ыa=ܨWT�민%i�Iy�H��
ɂ'=��J�hlC
��9e���W���8q#w�P��ysQ�R�Kv��d���i0�@7���^D�o~n�]�pC�E�Q#�d$_�6�L0��aP<�ǫR�Q��b���&�#hN`V6��۸֗��Q9P��x��ˀ�~uV��#�h6�eUIa-E��O�ʾ�ʮC�*;�O�X�)�4�������ٻ���T���_�	�)�4Ⱥ�3(+��Q�PA�K�&{�N�T�y!X�ˉoH%�$R�'���0<eȱ<��|��R5�(ʓ��8+�x8����^*��.#�&-cGi8W��+��F�����,x��gM�8:��>���"Em���2Mpҧ"`W��Nm,�g3�s��ß���b�`-O���!6ۭ�C����m�M�D/zN5"١c��r��5�1��P�SI?��l�nJ�D�*��F]9���*$��^4#�w�	����(��|w.;HHq���'�!t�O߾��`�y�'^QAS��}�[�e���t�NP����%��a{-h]�e�R�2�? �� �;��lpqq�Z�� �R#���|[�#�	�I}��1�߃{��/�r�<Nn�B��
�l���
-_`�)Z4X���q���J�[�)z����6�;��ߌWq.~@�+�|Ѥ����g�ML����Nt�h3��w/���@��(���@�f!��Y�a6������p#���Qm�q��/c�ʃ��.�LG$��+p������g�����[�8�h�?�K)��3[~�fA�����F���:OAj2fm�0Z�ú;ꈞ#x��G�{����&�:1�<�O���1SjQ�+$������f�CT��ʣ����nPK'��d�<�I,׆�R"��v@��Au����##i�?gQ����-z�<diz��! �B�h��h�c:���IG#1D��o{�4����3��1�-����[ۢ"�Rj�2k��{&�g��>u�4�<�^��h��fg�E�#Np�X��h���UV��>�����x���\/����l�C�)1�Ј#O۾\Z�z/�Zb݅q�G��+�%�C�c���@�]W�^-�1��:c��ڸ���;k���k�m'�3�9�kϠsp�*��oU��|�z��"��l^#�e������u�##�Yn4�dI�J���J��!���'�0.���LpH'�µ�֪�n��^���rݧ{͋9�'�]"��'x����\�&��.��tV�:-0��%� <�0��M/��9�WQG��FjK�M���Z�������w�I�ڜ�	����S{��g�pB	
�Ý���
NdG;�IaL���ԫ�[T�gd����S׍h���]�"��Q%�f)S��ۗcU#�/A.z�]E���VoX�L�u���F�`�PwQ�LKX]�l $�ۊ���a��fJ����t�5<t�l��1�����p���7�b�b����O�d���&TY��7�i=l	�����*fV�	�S@�k7Ua�L������?,�k�}S��FTo�O�8�����7�U§��iZU��V
(��yб����L���o#�H�i��&0�-�"~~>�Ě�x�`�V����{R��
�������1��Ҥ�3f��]泸.�n��=�ZL����ȯ�:�65�H�Y���c{/�z�?��J<^0��4���Yc�$+��9�=9�ۦUn��`4i=�dN�f�D$��	�2<͏��{ EAM��5��� �3�ǆ��I���:;N�Č��C�*D�@N�{�����9�$�aޒ�.�+_j:���4PK���"9G綞��k(>�W�e��ҟkp1�D���BH�d+����`���F�_%��aB��
���o_$B��Д҉Qo�r;}{��G+��ۨG^����%�^p@����D��O�i�=�����ȏg��hB�ǢG��k}�P��#���z�B���P<���9��w�2�R�2�� �!,��Azq�q����0��8]��-d���f�N:,]�#��kKY���� Y��@,�<��B<kմ��pH�}
��
�}�&��J�ٍ���Q�\ާ\�lГ����;��'"� ޴�o���~e9#���8�SE'�;v�+����b{�"%����Y]&J&���r�w��I�/<�T��F�܆]%��S�����(@�1�0���O�`�T�wM�ѽR��sO�<��(_,�+�*��L�IR!�t#{d�'t��A�X�=&m�a��%�Kn�B�����Ʒg�+p���at7́.���g8ER�����䞫c���UqV����9������{�eu���{����}������\��SA$aR`.ϛ{�p��C]xK޲�2������Zr��ܫj_��i)}�����G@zvO�#V�ʿ��V�m{���0��)�T{�Pr��D�j	i������� ��sW��b���Ǳ�����(���tw�s�g��Z��֒���&��Y3R6�~VE��K�PO,aə��X׸y�L[K�
��z���E�A�)��:	�@[��¤�En�xj!\�g�� �J>Q�#Z�1D4��:����O!O!lu��_7Sku�s�� �$-7� �Ka�G���|L���E��2��3��0/ ��6ٱa������{lS0�\ ����\�a�gt�T%��,\�S#vo�2�������� �zZJ��0 �����t��t���J^S�p�2��[F0~Q�d�%�E��F�� �ԒX�H���n��eP��v�Q��O�3�M�0��k0�j�C�%Ų��"E�Y1T0�|��-%8�!S@UQ���dĀY+)����Io7l��N%��}�;~5-�c�U��8o�i�U�U����ٳ˨�EܝX���^Xˋ'�*�qƮc����褢ɻ��~���h��{�3�}'������.;�p���XP��� �%&ҳi~�8�f.BC�w�
F�����x�%EXVmgWk���I�/�n��vI��SQ�с�y��p��t{���㾦��x�q��4��i�Ӥ���d?���;�;��ys!�s�V��G=<�Da@�
"�c�\"]�r�̬��6$X�]��J�фTT��pP��;��m�>�8V8s%F�mR��{��H�zo�@�;:�{D�w]�H�|�F��4Ur�G�d��X~���,�����H���t���g���ֲp�E��S���m��E�zF~��j%�$�E�uJLl�|`�
���({��\��&��t%�C�Q�?X͠L��*d�2`˧����YI����<�W<m���X��(�Xi�}A�b��	t(��Kl:�1G/eR;��d�DOlxMt
A2��ʏ3��b|(բ���;�c���cJ�O^qul��.��&`]E�f� F.؎3�i��ԓT�"��1@1����B� L=��k�s}��w���r��l��e���*�A}f��Z
�E��4�S��������W�`߈%r�̉O�}�=�2�'�od�3��$4���$~��H�:���-�3��c��h�V�@�������^�[��sJ;�
���u�ы�ѣ�>{�� ǷO6�g5�'w����d��\1
�|#�SջtqM�����$��̒%�r3��"�^�E����+�7t���j��A8C>�'dQ�
�s�e�E:��58�gx�8�~���в�>ؔe�ڭS�¶��
�>^�,�^a{�zԙ(s0C.h�Y�N$�D�	��_^��ZQ�����m�'5
n�(���bV]�({}�-u�2��D
��b�>���ԩ�ѥ����C�G��� B��Yp����vr�}�ɯ�_'lUdD\R����΍��]NI@|�D�M��)�v�-j���/��q�b��]�t�~�[�k�6X_��3$a�l�K
����=fǈ��4����^�!>�i�jl��tʳ��D��v�[(����V��4�<$`���#*�� %}E�o��|T!s�b�"��d8S�t*��e��/�v��_��l ��gd9f,����Y�[}�:���6�9���0� ��ߦMx���"���é���М22�2�..�r��/�J�7�3]ESN�����b��m���-3�X��%�������/����#��C�g��r��	�b���u'�b�H��"�ĘF@�^NL�t�_c�6���Oڪ�Y��ujo���t�����nV��p�.�J��¤AG_Ov�g�u��l�@b�?�{���WdC�Z�@%J��}ղ;����9Z��ц��6���.F��qZ�2ud%�3����l�7i{�B�;���o�*��( ,�V�b�M����S���є�A���E �7`*�'�7u`�Yc��}"����}���ST�!B_�y5	�>�TӗĜ�oؐ�Ƀv��fj��ps!O������/rM���#^��&�d��ߛ' �c|�`�y�ƴ82��Xu�v憒!����4M+B���n�z%5+Fo���Nh��<��|�=������O��rDƇ�0�.��?��H~�%
`�/D��U��a�~0p3������4Z�c':ʛ$O@/��A�s!w�&z��d�FpC�ƾ�������oV)�wP&����Nޤ ���B�0����t�!#wWjJQ�9��sƎmB_ֳ�����Goy