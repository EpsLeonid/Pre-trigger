XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��F���)��DSLv�,��?��S��r� ^��_f���D�O�4x�> l��fה�yw��m+ע0zC�d��=EM���m�K�,dsfL�?ȳ��\J�!J��~�9Jo��ɠ�����5F�ߘSk4ΗcuIE��=_�ԩ��-4"��F'l4�_�-툎���l[_��K�vk{'���*�y���57�S������*��LM{2[���`Bփߍ$��We��൪�W�߲^ev��m��m��>%#�-��>���h��U��6�ېj	(����o�?7��Fka�`�=!��ߐav0�����u>���:Y�R&�tGɸw;7<W)X&�1��&[�%�CR*�9�֫X�vt.&���
Y������o��n�f���[b��R�V�����tfe�5ms>��pHvN��Z���л6�g/��^IY,~<�s���ש��EI��;��;�?�߼�X@v��B�4|�E*��B�F/��4�)L���^z�͗,7����Lˌ��h�5��nyr�����Q�˰�"�Nx1���]���xpH�J}����bS�9�汚��;o'��oM��Y��YY5ԣ���:�LMÇ�*c+ˠ[�'Z���D�dư��~��9u��J�35cz��]��u|Q�o���4l�sZ���R��\�8��Ҽ�0
8�N��KН��J�oM�&�j`��b��AB�k�P�n�7-��� �Ч*<ĺv.�vucٮZ��2�XlxVHYEB    118c     6d0a��i)wǹ8Ģ���qM)���ܬx�(}jy���C��g��NKQq���Ӡ���J�F�N�)��H��M�	���ĝУ��}VX��p�3���)��?.��|�]ak�m�HT�Y@6�ٰD�b�z9�n���-y"f�������r�23���z��Ǌ˫�*	�p�n�D|ؓ�K�h�"�=,D.C+@�+�?�����y]�[���2P��=	�����{�
���Ū�⠷H�x3˨�)��@*d��sh���ގ$.i����>���Y;9���T����%o=Dr|����=����s��.��m��O�"S���T`�bS�\�W:�)qy�+R'=$�EZO�s�
�\�'\йp$G<s'�K��gܸ/��a���x�:X݆'W��������M��B�ϻgT��~����.B��^N�fwir0��H`U�U��؈��bg⠜;Pq�9����������r,���39���oQ��%S�A��Δ�5�cO����Q�J:�%?���:ŬjC���<�� �F���B�~�ì���t��e���mmz=�߀~B��"lrǴ��C[`�28F�3���>٪�xX��K/kj�n�������ICU/��z}���n{g��+>���R�5>��Lܺ��D���l��3͟�Nv�MRΨ���������45U� ��J�J� W8;s�\TYd�����h�)����%�Q�z`y���~�;���FFR!��>ZUX�7��,�s��4�{p��]�:P<33�Wo�E4F?� ����߯�	v��]�,N����и��@9IQ*�Q��E+�U�#
.Q�P�;�ii���<t%��{iq��>�z�?O	�]���n�-�*��tv9V�%��<��sc1��}�NA3��0o�8�L8/]������77g�Z��S�.yH ��Eةn)M6�1t&�������j(o#��Ht�,���v�<�8���U硽r�
}����#���鎒3��0@�s�y�`��H�?iH�ڬ3�V��B���/Zn
Ty�ŀ;���N���<���IH�g*�ޡ��l^"'�t���Ԣvg�EU���iG4���g%q�hWV�t�d���/X���*��%S�m���%��3��^1�P��[hR���9*��k��>1L��BNg0���ï��J��&���/|��man@�Q.8��N���G&�%��y����p4W�͚�;6��6g��R89�>�{Dx��А��cw��eH�c
�G������|��)6�f|S���O�
��+�����H�̃E;y�Oq�"�U|��V��Q.���E�?��p+�w�;P��xH�[-l}΄��n��D�G����K
���-�:�յ!b�[=%��}�d�!�ϯ���	)�y��M�6z�F������^���B�+�\'�����|���� �o][J�6�^p�3_|��ÈP9�Wc��m��a֚������87����@V-�^%E��G�W{/�s�s>�,/��p_���`%�MKw�H� U��߼+�pG"����m�X-���y2�m�}\(�o�pEy~�r�Z�pu��F�B���=P�\̞��rl������I%�eM"��ʹѱdw���Vb�A���CZ��eh��(f�$��X!�FRՑ�s<&�l�앬r���M�G��������� S��j�K����d�S�����