XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"���J�5��u|k<��k-��&�@�2�vg^����w�>#uCᬥs���6Qla��N:	H��OS9��V�]e5&�c7��J�ۺ>o*p���;�4��ǡ�XðsS���l�� ���}�9x��μ�נBy���.��T�zw
�XF�t<]s)*��s��u�����n1�-�ځ��AP]���
�H�!C۳�Kp%��6\�1�}���g�UF�v��������`�������եU�"�x\0������WE�y�kx����Y�� �E��H�~��~g��a�eP'q�>��$�i�6�zI]���G��l����fM �F} �O�4�9����e~���ZvB��\}X��,�+�鶖�*\v�� G��˙r]��Y���$�vC1n�:C�Zl�#&.xP��S��q���cП����+)%kq�5���h�nN��Nx) <Pd���tta�8e���k�9$l�e��lV�!����f@m^�T���$G�����X��NP���|@�	Ie�I����l_�'�X6h�1v�F��ۀ���^<��mƀ���t���QY�pd���^fS�<��1�h�~Ewd����2l����[�l�۔�(�速�@L���2�)�1���L�O<�^�	�1������K���l��d��vš� ���&w+ Lթ(��`Ri�̿D/ i�p��7�I�y�6'���p�;���x��v�{��]����Ղu05{��[64I6!^�XlxVHYEB    2442     ab0���hr�q���#-w=��opZ�F��E���P�.{(���A�C)Ԫº�@����(�5��;�Ј& v��(ijXS��A"*�d�D8�ZĠ�e��`��x�2A���yr��F�Cx\$����l&hS�@�f�:�EW�A�����y �_f+VƹT>�Bt.ң<nR򞡻�5ޔ�%C�6�^H�g�.��#��'.g��N���t�f�r��s+��ds��Gi�x ���$S�O�p�q$�}�cTZ┸���3t^`TL�; (�<�ApsBL,�ג�7%�F��+�<U�8�&V�M�5��]���	Z���]�OŜ���rFnΐ�,8��*�z��9��2��}���*�㚍��@Zʲ9� 7;���B�������w;�Fk+�n��������#%��P��F�e�e�E�: �Xc7b�/���Z�p �m��ok����?W0�8�V��\K�%����ZtH~�į�ͬWG",l�fk]����G��+mvR�Sb��}pK�K��X��K�í���B�GT���4��h�V�ؖn"��;��ׂ��G7yHMCv�;�d��.O�a�Tg���pJ�o�u lv�cܪ�.o�I��$a��Η��9W�%ח��r�a�Џ���}Yn(�p_����ʘ�<��e�ҡz��-iX�Ν��[�KpQ�C�
�y����6�%�3X#&	h��\�8��mEe�s��yT��<h�_��<h���}};pW�����b�������I�V���nVݍ��5zn+�����VaՈ��CClH�����?��(�'��Y�X�r���reԀ~dݷ��[|��(����y�={]�����.����3�Tk�V��Cm�-��4:+��`�K(
Ym%}L���0"|Է���L(dmO����\�v0�Y!�S/�n_W:�ۘXY���I`W����|@|QP�(;c�3j���֨�Z�Q�*���ۗ��E�(�$i���^d�mVv��)��+Lؾ$+:Q�O,��TK3� ]�]�`��9�i��"Tc�O�n��t��7l¼v���AXuJ���@B1LVw^0��!4�/�QDV�{��iJra�W�}v���۴����m]vn��\_����{W�����}H���f�).G.'��cPG"t~}Թ���یЖ]׉�&� jg�2 &�;�J�mDX�c-k"6S�d��x����eh��.�t��њ�.Q�J�N�EO`��8�%�\Ru����l�6#�X=�+���&����>�;:[���coiD<_L�N�;KVC�������TMf�� �}�?#�zym�p������h͟��t����}A$D��h������U�P�9��紽�0`� P���㶺�!������:H���@�?�L��&n���3�C+-��R���j�|j�MY�27�eqD�@E���}^�҄�+g#�0���T~"Lځ��a��9S���n홬�D܎;ھ=������#�䐢͚U�=ӛ~ݵ��'�y��R�j�A��#4tɻ-�b�Xl�/����F͛4��)wel�>e#�[e�m�j�W@����z��?(�󻫪[��&�#�GvY1�B�ŲdY@��L��#,� x3�N��|�[�}�����=Y�Q�@���h���d�f�1�}%�?F_�A�~��<�b�uCQ��r���8��q��'$���M�݃e�2���Iϟ�HZR*����%̖����`�����O����^�GR"NQ���m������ŽӚ����&(^t�)*I��.=�ATF��d�0l�5nc&��q7��04��
����ʗS��ȱQ��� �+ې�6ji�*�	��a��k���s[��<m�L����H�ɗ��b0Je��.���J^�t��4��{��[�IG�4��ew6���Q��?S��T^U��R>w��BH�w� ��E��Kښ&�>��xT����r�ݨ��� Kb"#��e�y&�5��Ԑɻ��=�c%2���D{k��a�K��������n�<��_��M����Q�[:�ؽ��,����)��W�l��f*	c�E��c>eL����7O�/F�����s�o��<Q��|L|l�_�^�'= Hs�Q�]��4yVX���#�]tN�����#���f���Z��E��;NUm�b������o�u%zO�I� �ae�[�����M 6s������_�Y�PZL�]d�5_V��<��%ӂ���55�|{X�1�}s���5"�lN΁��8V��ɊZ!3!�Z��R���.M�Z4'֏�����'�'z�J�̢�xM/'�ֲhA�ʶ���
|Wq�`�jĨ8�&�<l� '|>\�L��t��T�DwCZ���S�}6pKQ��\1����p8i��b��mo�8�S��qUt%�
��ːk�t��җ�����!&+�gD�;"e���^���ڃf��<zF�T�ˢ*�Y�-<���#�]U��  �h�*�"�W��uƍ��1dy��Ґ?7}(���+��[�<��u����;������X���BR��Bp��Nk���Ч}��8�È�;����ˡ��8�8�-=�4Bۗt�G����eL� ԧ*�ߕ�֣��iZi1������M�)=��!�B|�@6 �Er:pR_r�Pt*�3�߰T�q#.$��1��H���P��e�P�< H�QW-��/x�hl�ER��$���� #�s|�g��