XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������g6���C��S��_�7��F��:piL�i^�L��/��לY���H��� ��{�־-p�u��m�_�� ��{1�>.�N��o�F����ɠ���Ȟ̓�����dJB1�#�C$��������P������.H�((������~x�A3�Pt.���OL�1�*���H���UM���-�;��UP�;�b)�|Ir��Q��<��-�ݪ,��J�G�O*^%a����Q�%��Q)h햰��o�jτ���jois;wb�nKo��/��,8z(�U�ջ�5���������kVֿٙpt�ZZ�wܾ3c픫V��Ŗ�U���U[m�qr���$�quE]�3�r�ZZ}��۟��~52���/�;�09=��),�꜕,�Nh�<E�>�,�T.���ψA>�ς�"�:%�7���'�x�j��D&�-[�<)MթWR5��7`Q]+�nM;i�o=����$¸���de2��Gd�Uw:�S�J`�ӄ�|�F���D�,���bJ��۶��=�`�0�?���|�l6
9�
�/U�a�x�v`��y��n�[�V_�mm�j��*i|_~Ppb���7C��M�@j?
s���$�r_�fv�����%=����V���VSl����$rގ��7�_�T� �S�j�<y��Z#�I��]??+�Y �1��9�<��:A�<9s��^},�Z�+@��5�u �/�j��Lޓ���s��93����B�ɑ���Sr��-�E��mTCXlxVHYEB     f8b     650qF.��Ka��s��E�1�O�y0�۞|44+Z��>��3a���*�����B�;�mv���!��d;�	�qϣl3�у��������m|D�f�G%L�~�&J��錿>�9gTcM�a͌+�'T.�q1�7�{/�!X�̺DK�]m����N�.L�F�ͩ���x>�;4>���4��w.�3S�Jn�'V�.���f�v�\@���'j�M�z�!����7ci7�
l���	\s��Խ�sI�k5�ۢ�*�X�j�^��w�i���UƠ��V��+X������g�RHpdW�䗲�?�u��cs��T�d�~s$HS[��}M���k��Q�8�z��O	��i���edxA��>&�x7.�[�r��c�+$����8�w$;oxTݏ�f�l�\D��J7�O�����zE����j��ԛ�;�b���zk:O��R��wkl���<1����&��=w~'��'�8���ڕ�����C���A���I�D�,KP&b�K^k��X:�aN�����c��Ѐ�Tn��Js(��pTx�w�`39���0�y�4q�dظ݊v�*� .+�\�馏1È$�9>�b�T ���W/r��-�$�Eޘ�6Y	��8тl��Ԩ���R.�Ջl�R+���n0�<��(m���!��=��
���m-B���xJ����*C|N2٭�ϋ����0���&۠����#�woF.��=��?�̧��uE�=/T�QN��f�3Ekv���Se� =9�t����Ku�8���O��;^���'c��x]�e��т��Sk�k��d>c���>�dZ�=4�nbxhcB�S��eR\[sپE}�P[����։M9�<ToTq��;0�4>�d9���FH�6�Q%��N�@�Q��O�t� ��5��b*&(V�\̈́0��]�����j
�����t{�
�h`R�z��Iu���"ܽPNe�^v
VĈ擩Q���*bTe��V|'���+�E����I�f@v��팦��7��_��������5;d�NC<uC�_����B�V��HHVW�e��/X�.����t�����q�*֫D9!�N8F2�����7y� �M�F3%8�q.�F��?�N�r�*�{�X�#���O�u0͒��Ǐ?+�N��y4�଱j<w�����X�[��Q�/TG�A�V/�|�tT��<Ft���T�4����`��4!C�B_�e
9�4t�'��x݇��^��!��b��W�)�`�'n���q��X�!�c?V-�3��&) 0&�-%�BS����pa�G�_MHbW��9yQ��[\t2Qb�d����oz�Z!X�%� �_��� �C��`���~��F���s3�h���
���S��q���3։=(`*y�ɵ��[�b`d�J!�g�p;�)�\)��f��ܹk $�J�u���)��C��j���䐔�+�#��Ȁ'U���,���j��}ֲnӨ��@d<������
�x\ fo|�VJ�Ձ�*��y�GX�wD�#�r��\�n�2�&�}ی�=$J��$#��jv��}4�rL��}m�C���=�~�`r