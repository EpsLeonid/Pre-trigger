XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��c�F�99C*��g/���k�WAǧ��ܞLN9>D�z��9�>j�6��/HQ�G�qU���Q�����7�h�jcx�<��)�U����$�^�98�\n��Y���e4s?W� �]��e!+W�<�{�LcK�
XR��9��1@Ylj�D�8��S�� ':�]H�/+��2���er���狐7c$����1�y��l�o�:�f��CaL�M��Ҩ�6B�u�P�̆Mg&��^�5��D���A�����k���vj����Ճin���!H`��ݫ�O8L;-������̪��=�#�x���Em+�_(�Wp�i���:��7��7Z^1N��r�<QK
����e��&�1��5�>H�ɉd�������d7F==@�rӳ�VH��)�8���'{)�6��]
��ȏ��]��F
�>\��y���I֥�଑�Ec�@��Q�[)1�{�?����VR��O����9)��]P���R�sj$hzc��T"��c�j��V�H��X+nZ�#�f:��c_}3*8}J^�p���ϭoHCutk�{�j�,����g��+��ؼ�c+ِL�ˮ`��m��w�"��]�A7��Sɳ/�#�ILe�����>`L����Y�M%wj��L��\C��yd���%��D��i��6zV�In�,(�D�%��w3�>Y�t`�#SH���qF�ʸ�HM$U`�a=��y^V����(x��r��U�*n�uc�LÚ'E�آ#@���FB��[�gT���ܱ�_���EXlxVHYEB    1111     710�*<�0���}tй��^s�[�(�A(�c���{R�V�scV
�*���* ��|���b�Y?���=��?#0q=gZ={E�;,>�Ρ�F�/��4鹤k�l��W�U i�P��d�<]8Ĝ��9�'=a0��$6n����XRu�8��We�$)~nVjf���
�����4VA�8������0�O{z.���o� ����A���hBl����1_w�F	��ǹ�$-��y+��C0��ɖॡ������g�.Q�������B�t�O���������O�4�i�L�7��Q'����lL�1�N���S<�*���@�1����>�4�a �f��"r&fū����0�SȤ��R�[bZ�.�Z�P�4���*���q*
�o�^���~b���r�Vƿ_,�Ѵ�M©�>Qm����sh��� �_��A����9�/��F ��>��f03��#K��q ʩ��jp�H�V��@6@IQ��Ov�$~sB�{�\/�Ia�����R�!�q���t���ez�O�SE���BsQ��$dl)�P��S2�%@�v�,�2��|@����9���)7R_�q����2�	�^7@)�,0L�'\��ͱt�
-�)ǵ�G��j�n������L�i�(*�_�η'��o��ᖭ��	�ҙ���# �E�"�%��ɥѻ�)��0q�+	�0wT�*`΃0�gC�~2�l}�=���
O	U�����i�%���3�ЬwF/|��Y"���բ�3GK�.�����y�����ŀ��6��ߧ:��Ym��̱�^�1���i)=�0!hT!K^6ȁ=���{��[�[T�0�ݴx�0����	��5�������c ������S,���ݾ��H� ��=C�#���]��xkN�~C�|	�P�%{`��w�ۑz�S��k��7��[��ay��"�%@r�9���[��?iޓ��Sɫ(I?��C�_ L�i�5�VB�K��W��F$���{�?��o�"�=��Q���� �(��( %�U�^���6���74�1䛮��D�n�N����=q0��â�+��Ku�Z%�F"����7�n���^�@q�*C��Ҭ�R�"���;Y�{ #���.{�.g���5��T�iֆ��ɀ�����)���[5r�iM����q����t�Np���r�-hE8A����
�)o%<��}u���@Ukk�vBzh�g��C�)b��b�2��I���6���0W�@�!Y|s�[�gb��Ɛd�h����0�O���D\��(�=��~>���*��<!.GP�3$�j�u̾�!�r�i�����w�����A��\���q�j����������1&��ؠi���Y�����1?�!����On� ��ΎN�\�.�G�>c�C'�h��c���w�O_�(s~�X(M6��!��It�E�%�1�Ó�d�Bi�������@z�	���%�����X
.rɹ֎�8�U���O��ã3�:�������L}�����T(O񙹚��Wx�(v�$���eM=�,=aeO�s?~_ |pW��{���So@N�͞�$�*m��8�����*Q�%�+
�Äч@X�@��t����)�ez��ϩl^����=ϕqL���ę�6؀m��(�%6_�bo�;kU�'
8��Kߨ�Ze�;գAB�|����u��_ѱ�~�����þ鮤��H�%�2ࢀ4
���|ػ���mુ_���A5_�qS���h_��&�wC�kK�D���	5��&;�B