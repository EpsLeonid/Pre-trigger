XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����^�������U��ɀ�����3�1�/�z.�_O��Ys�0C�kVC�S����Ll6��L��@
Ї���e��9�f�R��]�l#���}q���V?$�Q�[��MN�eP�G���r���Lv'�s6�epS0�&�9� �澩�&�����A���fJ� �;
��Q�q�� �Y�tǪa�V"��/ �R�i��\��⛼~�U�����ۣX�\��B�]���pƒ��+��=~�=5��W�΄�:�S��$��V̧Qk#@8�晷��K(KVh�SN%ݓ�ܭ�mk\:�ʢf�󭜅%�$]%�5	.�x��%����Ʋ������{�bֆ�b�+�c�����9�(� HU��5
 �;���̙�9z�� ��2�f ���7	�Z�����C�9��`���c��-�vF���� �=?�4�<�,)��qYnC:w�n+W@b&���_���k��x��j��������/g�0)�5v#�qP~�!lb�H"�Oa�Qqύ6����A���n%˲��J��=�41¢\b�����ibTpH�fpǜHM���7��RF/曒w�5���z��Z�]��HQ? \��!�6�ә��&���V]���s���i�}4�u�	$碊���/G3ɰD*_r<x����R�S}��N�G	����50'`^�M�k�����P�|��'�M����Hۣ�lfv2Z[�N�8.A���TW�J�B�YGOK_��:��}L�� ���XlxVHYEB    4564    1270=�Öu
 � m��d��������쩘\=�d]{���{��֊�n������C�8q�d�>�mCRv�u�����8s�=�Un�������~����{fs����C�t����ZU렻CJb8����;w�b%`�iGq�Xs���d:�A�j>�v�&��+,����v	���F�-<t�E��gy+���k!ѓ�T��/T3�`"���S鴦��]3�@ ���^��P�R����K��\��*Gw,y!D	IL��rX�d8�*���R$��Ö`�E�gyT,�~����p_�R[2�-���Z��yI{]T��`lK�bz�DQ�u3'�+���
�^u��z\����Ԭ@�82g,�<��(1m�@�:lS�Ҙ%DtA㹢 9�F��;�8���?@L���M/IY�w����h��4�cWa��ۏ�9�/��	?�	M��	
A�D$�Jv�dR�s����z���R)��2��e�k��Bp-lO�]�?�
�i\���2�N%*�d�Ȫ�>/��k�"�Q���>�B���o>K�������\��P�H؊S���	�b��Ix��F	��Z��%w�bɞ؟3ݝ�m_�N޷*���!E�2h�iX���k�&��x�q{Ϧ���\�x��@�p�)wH�pN��ʽx��Ci������#������Nj�����&���B"#�W�6{%��;����D��â���S����J�&,�
R�7"�	��أ���5	���0 �9?����=���vc�PRUL`-�`��J*����r����l;YsP4�?8����1�5��	-���o�����(��{���ip�p��~�����v~>QT���7��)�X�p��_X�9�G�uU�A�.Yӻ��0���@Z���l�D"	W.�,�I6�djkq���^z��U�|���J�FZ��9�6�۵���Q5='i=����~������"�_ȹ4��W��Q�Y~cS����W���S�h���,�?{N�O�wcMBpT��>��;�Rc�~�v���:�L�X���W�=z$L$��&�ZJ2�g�60ZH�O�6���$ ��~�+HL&=�Y�߄ˉq!c�~c���vG��m�R�ДCfa�g��|�����,g<c-�]�(��&��������B��P�'���oXC�*վ��U�|Ք�Fh���G`()yq/���d;\+G_u,�ˬU��+#E��{�*/�Ȅkm#yZ_ۓs���'|;m� `�U5
��&wl~�:NJ�8�0X%�׽��N�q�i�'`J<�\t�|���D���I���?���ҰEG�~;s#Qxcׅ.!6���b:��5�/��$�Z7�q8V"v#V(}��8
@Urs_ϻ�Pމ���� � d�w���sTm<-1[�3`OZ�+�찕���[��;
*���5(�h�S�L��Ol�?W���< t;��d�~��8� ��gŸ��E� #�� M�.f�d�Ify�[@��m����<���� ���H7�M��5�n@�/��\���S))�o+H��{ytA��i��q��6���!���F��Sʩ0d��%b��!{$�~�k� n��U�b��:[q��{�?�_J���ǲJMt�1��K~��D��������ˡ�{%`��A�	�Wn��M�
�����wn�q�KF��}^8���cK{t@��Ƶ��6x^�����@	�}�R�.~a]!7X���`�f��Ts����B(e��)�n�zɔ�����j4�'FKɚ�K��jz���gA�����a�a q1h�����廓���COn_/�\a����]�q�rI��i��{\.D/���0�/�1��[�1yDʜrף��(�P�m�Md��3�4E����J7~��y|��c܍y��:"k^PQ6����e%d��g=�,��u1|�S*)H���g8�Qg�D졷cY���R�! w�$��'�x��=}"p/���E�ܛ&�V��4�rt5�i��	N�����_H� 7�;�Ax�D��������=�X"C������g�t����ö$�*��u���C�8����9�t������[Z!:Qy�[��=3x��&K�-��}�N�Q�;N �E_=+}ue'^�97�;�!�9O�'M��laH\��'2S��c1�Yb���~^����:��8�����]��8�ئ�Q$��jV&%�B�J�5:��ҹ7�;L�tcg�����|�.k�:���cki�CܖΙ@	2:C���'e�Mgt���5Q�;���
�1��ߟ@���B	'�>+4�N�vk.ny��p"W._Y}xg�i��ƪuܺ��ϚoG����Z9fNI ��\(�7'�]���F-�������y�At_O����oU�1�]�;Hel�Z�B}�Pd�w(.��h��j��6�l�Ð�)g�8h�+!2��{~��z�kZ+L�r�!!�!s1g]�A
�����l��٤ �..�t��V�c,��˰�(c�*it4����6��LM��L��250/Ǡ��N�������Bŝ�X��
�̀��֨I܊G�-a߉����Vm#V����,'��Y&+�X0�Λ=���bE��O��D��'�xN�)Y�|�:�"}t%�M\��=a�G���9M�쨧L�n�~�P��V�H1�Kq�.�b�Z@�Q�jnNu���{�f�`�s=-�̞�X�;�w��)��"L�կ�� 9�6c��xb�ao��w��,!�^�E��h'��M�[c(��q�$&���R�+ܔ]
�3�juD�ߘ9`�so���*�2��[s�Cr����`�ǟ��$�"�޴�����x���b
�����]��jP� ��C=�l����>�j������Q��ju�0��������L��IAB�ң�h!����*mlO�RX�-�a!��@�}$.g��t�KBdH�b0#\d��x�UW-���G�����۫B���\���<���'�D��$t�����@�ꮮ4S��OD��C՛Y��C�UM�VC~�m/����. L�{���������z������24 4z�4��ЅP��Q?0V��7j��p0N�i�O���8	R���\3O"�I�68�47����0f�����bS�w�����Ux��&!3�z9�?s���	����D�g:h�ϩ$��H�j��{j2=a�ČE�Tb��dNι�Xp�H?�X�
?}悇v"�� ��C=��c*���h��)��E���#�uż����Km�$�X�i=R�J��U$��`쮬J��0eϱ񫋤j.Yv�w�c2m
�+B3}3Z�Ο̱6�_7�[��s����Ճ*� ӹU��a
n�����&��^Һ��&��^MU����K����2��=��UI��� ���h�ʡ����t���8.R\T�#�4)2�-^-�6:�F�*�uĠi]�́��HLSWv��-ϗaG� ��e&X���GS�
�����x�r��͇�Rp�1 �4���Md�B�����^)����6�6�����*�u;s�� ��0�B��T4���ɤ�A5\�~3�u��_\N(�sv����埆��2X&�;��W�~^8C�\��T���0�+��g������StX:u��^^�0�����U�V��w��c ��{F@v/��v�y�����HʖM��4��_d�n�HF�v��-�����{�㕀����,�ρԜ�΄���X����QV����V��B�X�0�-P�L/w"J�j��ް��&���@{�7ˀ�>Ny	~?Cz�gOSA�4���n�
0�u����U	���j�OCK=��'1;mϐn�4������+"#��P`Ĕ�놿�2��������?�J��M�*�5�6�Y-5'�qb��gþ:)�
.jz0�?��g�?q�m���e� /G�s=���G�%y-��>�������9��TP04�$�
�OI��b���ATF�TE.�-��ڴ��T�\�(�`���f]#��H��OZ�;�p.`����"@�TwrCp{p��"^QiDrSNEdό��u�yݡnZ���?�:�k-I\�riʺ�v����K�*,��4�����׃��
8��Rֈ~J �4���v�O�Ы7F��X�a8���U�3`���\��u�"�2�F��T@�|r�}��L�����˲/i��3�F�D��[b���Wv��GH��&R��3�{��������`!O0��-*&4�nE4�	A���}� ��WZ�<ơ.&8��ϖ��q���!d��K�}�����Ú}��p�Y� H�9�R���7��J0�aAo"��	��T�`�'d �E��ܐ;���W.݈�!\�'^iO3���#���șZ\�S��X6���5=��z�&�Z;�H�N��=�ec3+�ެ� 
$1R�dI�x�돯�^T�-Q�Ceĉ�N��\>�yt�pr!��v�U��f��Ao5X�)��stx^Y3��s1���}o��:���4s�����q%E�I((MY�f�6��d�%��_f���4m��3�@-����尬Cu��&P�d^��lv�9��`J7��˚�`�ގ�z	������r��n��B�I�������`BV��d��T��kM i��/�QC�w�.8�s�)Š���: