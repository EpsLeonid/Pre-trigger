XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������c�R-��'���j<6�6�*?�����xp�ȭ�����y�d�0Hј`O�p!�kX�p!BM�؀P��p�S��B�̀3^x���{X��Ύ�(�r?=Wg��x,��m?m��\~Sv���b��T�`Ev7K�,�:�Ǭw�����+7�|��8�j	0.@����Q!�rt��⟋��, u{v6�H�q�>�
q3*��,V.��}o�o]�.���!V��J�O�nP(�ly��ʠ��ߓ�쩯���}����Qv2�]��G�8v'�Y��pn#�l,�Eto\L,iؔ���W�|��` 6 䨷�3���$;�YF��H�t/3�m����q�n��l/�n{/� D��6����\e0.��,wwi��o:�� ��nB�e�iw -�"�'�Ю��K���8"�Sh�x|�d��]q��߀u��$�Pe��6Eą��[��>��Zj���b_�0��D��Ò���c�M�\U�f���gKq��śr'	87�F���r���l��M���\��g�_����T�M�P�jbfy��*�4�a�9�ِ�Z^V��Y��%*�l[�R#t�\�5x&c�� ��3٘`N���F��@�O�0���x9��b��L^WL���4$R���	`N�u��)4'W�ʝ܇g'BJQ��K��R���'.��P�,�ߜ��S=%�T[��xh$�����9�ӱgw�'0��M�/D�7���quj�$c�Xt�B���H�%�������C$p��XlxVHYEB    38a4     d00����B�KZt���_T�&cP�v�Ҕ�4$1S� wuHl~����-��u�$�{��I���p�Q�ź�
���pLi.��(�ّ(����i��ִU���o�c���.T/b�>Z�?r�af�?4i��s0,��q�%��,=�D|5bi#3-�#�ҩ�����i�-y�ku-�W6�ԷhO"x��4^��s�WIg��)�#���\�Um޹?���X�ÈV�a	. �����q'����뀏)ǲ߲�8^�����}��.����o��EB��x�8,J�̶�S���:�9�3��Y�Ȓ���#á�a�~Qk����+Gs�W�}�7�Uu����W!J�^��Kp�#:V����g}�6�Kv�/ڵ���~*ł���,��$�Na g
_8ONLf�\�#�.A�������������r���Źя�]��%��u��W�: Ώ��9����W��%N��m�,
n~��=:
�O�7�Г�+�\�v�g��@~�,T�e�a�43���)��:�8M&�o;n������njL�<��{�{7��V(�hQ|�!o_�Q)��bT2�,�(���, ����d�|{�*,u��_l��FX���RT�ZEt\6��D���ׅ��iՏ���'�fy91��{xD�OsʸU�������$����p���$S����ص�x�b0�L�wb�`�
#�&��Fnf7���E�#��S�%�j0^:nFU��_C���o-;<00=�Ɲ���#.G �WbN��=��Ʉ',�	��q��gh��,�j��&��R�U�1λ1�
�u���,CH�c��/4ᙁI1�NĞ|�,pϻ�}�7u׃a��R����p��i��RCl>G/�(�	Q#��@NY���(�u����w�x"��9$��N�OR��_44s�8�PDAt�@�8ZZ�cp� �$zu<������N=�?�;���0��z�	�Υ4��%���P�Y+�?�>ʦ|n^�_P0��H������_t����$$aCBV������R���gL�_"����#A�պж9�O�b�r!5,o�lPLޏ�s=�UE�Lwz�:/��:^�}ZO��1���1���p�,}��y&�sZT��,�`:#||��?�x�����S����3=FF!��R��:kJ�ޤ?�4�L��^��e!���eX3�E��M�,����S�9�㛢�z�_:ζ5���A�)����#T�DDLM',!�w��k�6�q��}
 �Z��3�2׷]'D����RD6�1�Q�]��F�=O�/p�w��aN^M�2Pel���{~&������P8�9.|�0�*)b���Xb*m{ŞR"|D�V�������x��(B���C��+�por�;�2���x�����Y���}��<70��"�o7$�2xxq ۔|��n���k��%o�ߛ:2N)[�K�[�8F�"4g�f�Bͼ��V�|��S���In���ܺO�p�ls*��]S�G�e��z�d8�,���\���x�w�r�a�F���h�2S�A����G�It�݌ᖱ<��r
~l:��,�����mkp��UkA"��6#E���~~�(0e�1��*	��A4g�0,�?D�< �D�"�B��r��R�Y��%�f�TA���nj�vPŎ�9�+�<��7q�Ar�3t4�M�h��W�R��a�p_��R���NrZ��I���0
�7t|*����#�����4.�;8.$�k(�}���$�sھ�3�K0����<<K���F]p���1VPF?݅o w�纃�$���,��ד72F�uܝ?�+E?"�Ќ|��r�#~�!M<�������\�3儁�5MK�h/��(��s���g��<�t~�h�(��1x���߼�w����L�} ��`��k�!6�,'Z%��bvX�4��h�zI���I�	�������>�X�'
~Q��r,�$��!d�Q�Npg����,�|���<��A���9
��L�2�&yx���ޮ�� �UF.����(�&r�����k6И�����3�?aX2!l��JV�2)-����hp��צ�qJ����I_J��Cq��a$,T|C���G���j���_M�W��$����"��t_��:�<�3r�:��ox���#�7�Ф�3;�N�����ö��x*�	�=����G�F�BB^!c��)��M.�ۜ��Y����%<��qC�ߏIА�V����|�rS%,19\��OB7�}c��	Ӳ��u�k���I��J*6DWZyR�����U���)o�,����ç� ���Q~d�N8=��U4��Y���'�x��'��tΤ8��n$nJFu@�49=;�������N��y�b�����y3����*�D�6�5EL)��z��k�¿x�`�/�`|)��8�xQ��`Dy� �>j�É�HE�
@½���IƵ��L� r���'U���׹�-0�'�P�-m�g�r�ؿ�vƦ�,vcA�}
ߙ��Yw?�Ju��
��-K�5L~�.�)5�OĘ�cu��!�`�+��aZ����6^d7����i,L��h�+)�Q7�B��L�Q��"C���i3誙��/��B!��6���e�Y,�Jj�	����GQ��Mz�	��Z8EC%������J;^�:�SWo3ǩ��"dA��&`�nF�!$�o���ÿ����h��k��:�(l���qdl�O��DQ����k�6}&7��?�+��#x���?LvxaO�N5D��%���az�F�SYc�-FP6=6��_�S_�c@�0��!�me5ˊ�rƟM~B
a'P����_�5rS�r�c_�z|Q�D��-@��ee�R?�������p���2���8'+�~����W �"m*,�<�M[v�=�{|,�[=P��x�t��4�5�d���m��l҃9jq�,��u�sg�O�/X�4;l��T�5�4��j�H̑74I"*'E��8t�?�A�g�Oו��~��e�V{�D�������q�CE��DlM�ww�Y�8���-=�<u%A�"��Ol(�=j׫}F��XZ�ur���D~��DbV^�Z`]���.'-��b��Bf��!���N���3�^"_Lc@����7=�@K�ų�t���S1���1�uCA�j�����),�T��3�$� y�j�gZaaH�Ѥ����dj�*fSaS��Zk@<s�|��Qk%�qP]�Վe�
fQ�Rqp��0@*Ʉ�ͬ�5��5gWnP�^�ފa:'��