XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����A�? P7�j��_�(�S"��={�#
����-L�|�����¢;q����iM|`�������T���ve�;̜t/�Ûu�Ź���e�%!良>���"˂5���Qk�I����" �1��M�1�@'�b��z@{�/��ài�U.B� ����b	BPe�(�⨾Bm�����	0����FX��3�+�2*'A�~	�Һ&׉ɤ���p� �N�^T!v_g���ū=k
����t�P�m�n[���D��v�R�m���5ܝV�`�q\��n�zvn�<��=`J��ѯ/�x/r���ȼ N�bB��e��ؑy�]��AQ��^4���$�����FV&)i���lN&:GH���>�<�z��nT���ib�h��D�)>�o��Q"*>�D�iX�����@q�h�`+�@
�(Yi|m�8M_���L�T6x�mz*۾����!��Z|b^m�0��`~U��c���OCtsJp�� ���|�
/�t֝"Q��v��ۿ"a��Ŏg���F�#�F�67xWy�K�)����X�+��ZY"�އ�1&^""/ާ]̾I�t{<�� �6������:�)�h�U����(����#F�g�#���#D6Z�ʒ&`gY���2^��~�琦��F�����9'S�BמBQ��ٺWl7�~�F�G�bu`����:��jѐuP?��?����6���e�R����:a���J\	%Jg���?93gE�˺)T�1�~�����&͍����l9����XlxVHYEB    9653    1860�>7s��?T?u��uU��˘_���!�z��ʰ̴ew�bZ��&�v��q�B�xP
���F�{�x��\���zɽ�#�����$Q��}�tT�Ý{�"����96$]�ᬫ�;�f�.�Ğv3�H��'�~���8�6�a���:e*�KA�z����;�"�1w|�3#[��2u��F_��\сД���#9k�όiM�%{t�y�)z�_����ݴ��x�%2��2���?��_�����/>n���e<����O�6n#���z�}��j#�Ǆ�0܆M��n��c�e�Blx�.����6��s�2!}�O(H��_�o?hѨ�[: ��u�y��4�ad��8|�@8W�?�k�k�|wӨ�u�'d/���2Eߦ�����Pc�Y
8H��|g���~�V�6=���؎�H#�~s��K&�M�rP޵az!|��9���ޟ��ir���^T��4�+�C^�R; Ɛp蜗���������-�V~����?�5qm|Є��u��ʂ܄�N�3�7��w��^$d����A��ώ��o�7*Mu8���W�3���NȄ�
vz�1���}	�M�@��:<=������&m~v+F�scu�������.�-,MJ�e��� u���yD�+܁S4Y�ـ�u������\�ѸޢV	��T\@��H&��H��+���N�m�vS�����,�å��=Ѫ�4��Y�`,�H�%�ލ�I�Q�#�ο� � '��h�D�0ub������d��ڵW=�R�LDgY���Q��{"HA@E�n�ѸU�$�k7�)�ai�w����E�A�=X�䱓u>��m�|�-��Q���<T�g$��8?�:��W ������ɥ���i����M ���X�'a�f)�����CTA���{A=K\����SlL_���:��(L�������Vu~E]:Yi�|�q=7�4��)��WX�iT_F�&�I�C����2�z��R�ۢ�Nw�{�<וDq@?O�ɋo�	$�g</�[U%���E�Cĝ���Eb�R���g�Ҹű�\��#yp�����s�����\Mt���g�"�y"Ğ�:M�n��FNZG������yԮR
��DΆB�/�TԹm�-ΚS���-'��U5$��&�ڗ��OV�<ZF�fb�so��9�.(,�}33�g�zr��8��DA+ F�n<�
Sߎ?�
��eS:������D΁f,��I�����7�:�`�_>PU�q� !%�����3�p���i�$r���h�)Mq_ި��lV�q<�`��_��� �ؙO��jJ��Ci�a %��K�n�Đo����-U�X�3R(�5�ݹ�7�dĥ��d ��7?܌����c�.��th���/���Ǘ�ļ��Q��'���#>��^�4��es�J�U����̏�#�J��޿��rMUa�hip�G����٥��/�����k��Y�j�}#�e�ZAi��Z
��k7��6�v��Ӭ���b B�~�u�ӛH�!����xk9�
�y��aW>Ӆ�o�����ǹ��y-�4kcB�я×4��!و[�z��ʙ�,��Ⱥ��T�o��h����<�xd�Q��p�@��	7�8t:�Vߣe��T� `�&���N��U���/sS���5r1P�3OM|��6n�@�zG΅�yP#m'���	d�8W���3szn�_���|��(�YY���=4���=�5�k2�A"h�4]V#��.m��(�^����M��n�џ��h��� {��*|��_�J�4�����\c"�����֘f$�C��|�d'�۵O�礡ս�rk�\�7�=@����-5Oz �]HJC`��z�M�&�t��ҋ�;��^Qrp�0W��YU�w��J+CLl��]��R �-���Z~�mcHF���!�����bӏ����&��\+7���_��h��_�%�g:���L���騺�\�P��h� ���F�`q�8L2#~�*Ph|{���>��\|Ⱥ+��]W.��)�&��̖���=�eg�Z�@I��#1�L��צ�b��H/c�ʀ�ݔ����Iz:�T�f����~� �6�Ob���3S��;��2�d{�AieO������iEŀ[Dp�.�W~*o��y��>6%��ӎ��˸B��_�vV�}��L9�ƈ)��3�D7X;�ztEC�����W����;:���)�@�)�dp�̫���y��z��Cd�m�J�f�d�V��y��7�)=�P�{�w����)J29���M�!6�J�����h^�xߥ��hIX�l���C��%|���S>��	N�p�Q��@O��?B��S2c��+��(�]�1�y��UƗ��ʩI��|eIg�H������.���*��r��, ������������
��\���ۮ�'\�����ʶ�^+J+*C��8��Ҙ�G0ӡ��:�̄pA����7����H%챎��; �>��t��
��D�%�ئݒ�fCx�J�0��,����4��<��P��������E%��̽P/��	M��9����D׭�q�t�L�g��(V��0$R������ s�����9g�Ƥ�$��L����W��EX	��v�,.�*J��.aJ.>b�ck��S��P��y U�[RSp/,kũ�S�<E\���yR �7''���|�"G����^4ɫ���V��:
e��D��DuR�x�##�!ի�ݵG�fe��؃��ע��&w���P��f���!�p{��~�� x|G�3(��S�� ����\�N��� ���Hhz"*�|T�a)&~�推܋�E;�h�@^�V��N�/�=سoLՖ����kQM��� WV�����	�wx�X^��R��"�Hԑx�mSxlU
R����)�HH�6�9KH��mԞ����Ȭ�އ��/,�ϫ�͘|��Кƪ��4��ß=v~�'�3M֛�#��D��CU�tUOI%��E��YӃ�4��n�
�`�1����H{e��U������Vq�ǌ�y �5���	_�l,�"��T���j���"4��a�P"$��d�}e𱱜{�	O�W�skP��pu|���5�3k���V,�[�L�i�(�l�cl3#�����q����ѻ�>��lˀ'M)����?�j~o�o�9p<,(J[x6�,�s����Ry{~�eѝ��\��1T��jo��[����J�Q��~�����k&1#s�D�������x2�v��R���v�������h����h��ZF��_���*�T��iբ�i��=`XK�ዽ�;�d3C��@-�J�N�܆���o�y�(2�I��II�=i׹�m�Rv��c�S�Rʄ�J��o�ElvK�Z�+��/2����v!��P#��l���v���=�Ll/A��>�
R|�mU������'���V�D�C���^7be����'J�,y�dN�ⶮ|��q�������Xo4�L�UA�7~7��m߉�sA����o�no��W�P�k��|��w(�(�>�W 6�$���Wv���yfa[t�B����_������i�{#A4�O�R�,zA��}���Q�3F��,7��x";��t����4�P����v�U�����$��;�jrR��~�T�,��1t�!�<k�t�������aD�w;g5+������0"����ȃ��'Z�U��H��,`��V�{ �6W����'���3CA���D��6������衯�gE��ӱ��.��.��"u�T�ȴB<16�}���% �sno|�B-�6�}�(��ݠ��a��@�V���`x��JL���7-h�ܩZ&�o���{��#�pT�j��|(]ɂId������z�C�� `y�����"���Q��iH�	�� )��'=��� :iE�In�3�;��D���	/{��c�W��'�� w����5�,�@�v'XQo#S\T���E����q�'m�+[B�0Y���&���W��s_�"t�6"�6Y�2ӣ���H�(s�5�������
o\L#�յ3���3$�&i���).��~�c��٬w�ZP]�?�^#s޹�m%�����t^��0� ��s�v����I-����yĐ��������[y^���O��Z0�A�Ωl�:	�p�ܩxf��^X���U� �F�|
;]�_�M-�Q�Q���a��G̵�@W����$5%���_4ߦ���x= A
��R�8�tM�Hs�DW,^({e@t��J.�g�>����D�+�uW4Y���b9ZW.����=n�����!��%���~߅,���g8I��s�����])P�!:�{��m�+s�4���B��+�:,��71/��S�vew61��?KՉ��%˵���쒙 Y����"��qA������3�ec��mGp9��Ȓ�N��u�����6K�Ab��/E�e<,R8qȩ�H_X!$z�Wȸ*F؍ԟ<~3v��ō`jM�3��]�q���)�<H��Ϲd�Gj�ϸQ�:�����,�!	���#�p�8���(��������*�A ���X�+��Y��\ޒ�D�=n%:�;�MF?��wM+:ʊX�s`���xfJм�F��f1&�щ�ߢR��5��T�3d=S-�N�ޙ��KL��y�U>�E�C��P3>�vz����*U�Ӊ��KŎ.;��$��{�S�NFj��kH��N�a�NW�֥yb�dI�������+,�m�j�:�!�]d>=��r����uŤb୶c���d�(v�ܚ�ڏ��2J<؛��'�r0���wz2gh����o�R��(}��S�/5~ﻑ����d��=|G���%�����ps_������W�g��^�<�Qa�Z�W4zJ�3�ẘ-=�s��a����?�P���_Ь�]t��G&PJ�^;@|�����"�*N�8����j��&$��`�8���[�
N��-Ǟ�Q�y�&Ef۫e�88pv2���ג�	G���:9:5~���>�B����f���:;x'��M�<Vϛ��~q�e��q�7�O�Z�kA[.EM6O�V��R�m�'R�ot �L�s�D��͘x?Y����:�[~H�P�W)��5Zl�wF�X�K⚐�m+�!�/�c�l�k�Ӽr���3XRGZMc~4�bEA���q,'�	1i�^~D��\#������'��e:B��T�T�2h��J���o_���f�	�k�:~�&
hwE���˷z`c�OY��,d������I�sA�G���",Q��_��Ȅ��V����Ԏ��r���7s:C��>�w�æ������2U�3%���3" ��-�j�/-MH��ll������#��D��jW�8�<�A>�L�������O1�4�#��J�����(X=0�^.����6����i6_�i���b�TY�K�ZD t��q�.����!W�B�� _C$��1'y��wd�1����<g��t�i��m3��*j�@.��K�o�5���{�#����gp�~]�"�s��B�/(�DG�+��=�QN���T�ƞ��U-�hDbQ����������T������*P�'Z�+E�[�.��.��˯�m#'� `b�%�5[X郎��NY�w(yX;*�
�X:���n�йl���pq^������`?��u�{�4�cl;�usy��
��3�����c>WW����6D+�x��=�t�{;����/�?�T�c3:Պ*�ǻ�A�%�
2hj5l�Np?���ؿ��$H�R�d��߬9�&���$���"��9��0�n"��y��l�����-k���j�.#%
5�u�#����$:S=%BĔRLuAOw[r���%��:f��z�˲�f@1A8�(�����n�f�EA�UN~�1��>o`�Ngmo��]�}+_b*�}r1��]�81��'^�R�V�;(�[;���˝V:���ٳAHe .߷n�v�6c�[��g[��}�Y�Dt��p��H�WĪ�tM�@A�*����i4ۛǗ��	���&�Ž�x��E)�SK��x�Ĉs:`�%`��$�j��X����{L��B�暴���(���u���9�����~�b�t���&�x�^�,�8N��'�8