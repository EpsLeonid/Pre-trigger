XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z�=E��9>�S\�N��ħg;C�iis~d�6�S8�'��G��_a�0��T[�[W���"*�bI�'��D/�Z�v!z�Y<|[�"��e��Z�gx!M�KS��EN䦹b7 {�Â-�Z���z��\.\Gռ��~��:���~;�_OVG9)~>E��+����FK���< ���h\�z�dV��d;,ʍ�����4HX2Q)��D	�!TB+k��7#�*�[J��#K��*C�G����O*�{Z�
U�@��q�i��@R6�w#j�5��^�d	�
�2W:�Q ڳ(��l1:�e�����2�I�d�ǒƭ~d��<Z�(j���2��.�eW�W�B5c?�D+��;��s������I{�;$H��i�&�sÀ`MP6��tn�P%<C����<y�
�#����=����{��*o#3�#+�xƀ�[L\�e�z1]/���_h$��"8����Ƶ.d��8星4j`g��i�%^;��C�5)G��櫹-@��9�]b�"O��a���T�+ a7¨�6��Bk��X#��&g�_р��V⹙����c�iJ&�!��}.��$����w蒡���m�5PM�EUg����S`x"�J�Fam ���u��è�C�i娒[�öl��ive�z��J�:N�0h'/�?vB1��ɰDM��h�h�5^�A�t*��b���Ԩʂ���"�\4dX���-mW«�i�g��t.���v���U�	���ƻX��R}��a��9��ڿ3GF	udJ~V�XlxVHYEB    4564    1270|�B�ح�'�k�N����o�m%��p��#����_\��QNa�,�~5�{C��(�E�0Q��ڑ
��ٱЀѷS6��_�F^�80�q܃�K��l��GN�I.�tm����X��bF��+$����!�y���6�M��i�ř򆇫�'���ʢ������h�KJ�	��|6���jf�>˧��x������AjNwHځ�\����m��s/= �����J�^76p��W�VD
�x��C:��V�U=X�?K
&��I�H>�=:�̤T��"��{����}��t��.MG܉�A!I���%snP���Z}6�ޮ�X�ȋT������{����k1,�|���cAz$����͚��rij���K1��sܳ�vti�y���ۦm��?@�.V��sZ`�?%I���	'�����đw_9�kB�[dƕ��u��O�5��?�\��XZ����!K{�;u�nO�۷�b�Lq�Ó��z5���I�����'�w�B'���#�</\F"�]gD��)���k\�k�i��q�<�:s��xn|�#
��9D����A�	r.��xն�~�/�Ȼ�A�i��U�pTm���[N�ReF[�v5�c鄭=j�~��lRi$2�1����g&��R���Pn"�P| ��N6n~Z����sU�u�YI����h>ŮP����7u�!i&~���d��8g��MY�\�c�!�W���u��������S�R�>�SLV��ʹ��Bo���M�R���CF�PD�KP��
6�P�W:�j���ܨ��◯��m�R&F��%S=� PB�sM�dF�W�qK�����9�W����-Bq��./?@|Gh�qϭ/22�|n��>�'�L�5��/��rq}VÓ\h���.�eE
���"B���.�Y�Z�Cع���6���z�����]Ϸ�	��s7�Y3���ȼ�3�	ɩ�����A���&��M􎹶��ő٘d�x����i��㰲ƻ2-o�~~�j;��xF�C ���1�+D����,!�J���<��T�.+��c�5

ṧ]����g�6w0׳�-���R=�b����c�^4aE��9���� XY��Rܔ@�����|J��{^��k��ݿk4s/��.�1ư��~��{�/)�W��wJ+/ֽ��]P�$ԪoWh�7�.� �֕@+�;��Li݋� ]����J�6�(��W�p7�"9(�E��-�d9�M���.w+���Dӳ;���|�3�o��e/�q�眰c�ԅT�
���Jh��e�N�k���Bh^���
�gZn�\;�0J��_�\��.4Jه#��/գ⇽�&#|�9���z҄��F ��L��,����b#�,�q�2�o�9Y����D����CZ75�+�����$����&+��I)�'�YH	�~��
&ڰ�3%�/Ȫx\-�a]\�=>��5--�2C���#ֹ�������;&&3"c�YЬL�_~IV�'VQE��C-��~I�!��Txַ�+n�x��c�U�M��(�/���%\�4ܻ�(��ž"ՈLM���K7�X4\��0�I����"�<�^��S�v�;Bq�&�W���@9�1�C�ۉ��������Y�/t�p6�<���v�&���D��ف)N�l]����Eᵧ�(�G���B��h��4բ�����tM�}1�Ԯ�0��i�x9�A��A\DTZ�ꫵUn}Fl�� R�evs@������+�TU�k��:UO�����Ô�3�6�L&-*k�X�'�j#�ڦ
ϳsǳ�F��gG8����n��g9����p��Ó!/�X@�p5�to36�ۭ��;�<��5J�Nj���~',����ȡ�Rc�����{aN�F��*Jm!�J�0����
%�\��1�Mb�R��	B.ϧl'�Rj��En�w�*6+�o/��3��ũ� ��l��0dh4�
�E��Gr��t<�\������k ��v�i�����A�.f�at⍌�}�� �er�5��MZR;���TK���$���k
A�O�+����д���(�胕�L�������R�i�_.��uxtڒ�2 '���*�*|L��%��2�b�e�����`��9��?�&��#z��&�(c�o���q���*v�ٟ dQ>(<{0�P� �wx2�P��'�2�-�ģ�8�`�M��T��3��@�����_N�־�����"�zί+�v;w\�\���+�+����*�0b�+�LFTϽۯt+�"�8[йib���T�wH�*�j��9N�O� �Ab�qq�)�!����]���YCa����3�z��!��W��.��:mO��,b��
��L�� �E`ίFQYE
si5Нr�-8�~H6��<H�,��#D�H�㇑@#&,#�×�
۬a��r�@.��D�C���M�����}�F�
'������J̴�,x��:�p�z	^�fP�!9��gV�P��|	�P������,Md�}ͅ)��ae���M��%(��|�H~cH���+�i��lZ4~A�� ���Ǝ�(�v���q�͵�s�a�Pz"�
>8^bwE�����\x����Kn5��<��1H�	V�� ܫ�NK�j����
�Z�+����O�F�G����6��~9�2~��w����L:��(��jD�;I�D��s�B?$��i�wr:��`,Hv-��PyhzҖ"��IX�� �f������RD��χ�R�T�_ ��+��	4&dS�z�p4�2ȭE[&c�<��)��"�����n8a�B�h�{ML�
]����v��
�θ���f�,�M#y�/�2�uo�"G.�=�2�l7	�bj�U)�>��9��ɓSN	��Q������_U�þ#�_�h��ۓfJ��8�~դ�+��=&��7�5�"��*�3cU�RPe�X�� �le�?���QYF���.���}���mƣ.TT'��3+�F��d���d����b�����,��������ʦ	�}�����뚄�[B�C�\0hYd:xze��4��k��{��+�_�X^	����s Xw�i-�M=�0\�`��o_�7�i��G��)�޹���i��[ f:Ȇ�;�F�J�d�Ng�	{��v�­�Q�{��Y��˂��۸\�-ݳ�O��M�r({z�u�}1IpHʸ�!�g�E6�;�7M�eV}��oZ�����[j�$C�*�@4�ԓp�Jo�Ha���T�Lc���?2Rn�?�i�k�/�*ڌyB�zLf�)�0��ԏ���&���qa�o�=���<=:2�����"L��/q�G�>�$+!��#�Y��&G�����{-I�/���y�V���CS�DZ����<�ؒg���/68�d�q���iVR��I'|[M��\Le�!<���'wg��}��܅�?�Ԧԍ5�3>5��N3Mm�
9�^;�K�e���[t�m�^����ҏ!���§�Y@�SHD:O�����z�U��ϡ�i����:l���V5�;[���)b!b�G��b�(
��<`a��Ӝ����D�O�s�m���8`1yq��9%�'�q���%*�U�@B��:ak�srUU�pݗ1������ٜ�h�I/V@�r��U�6�˅���|����W"���Ӈͨk��"�fxi.T��(21q'�q���n������]q��eJ٣�{�1���>����!ؽ{h���/׹XJ��^�G!� ��>�����"e�Ƣw�}PX�X�7�y�W���#wTA����_��1'�Q�ٙư�L}��wW(��y2�N	~�����9 
�sg����wТ9��������S��b�hD��z�%,�b��R�fubȈ+[B%h��� ���[��c��p��<a�O���Kp"�yB������,��E�� yi�!/��sv�-%�Ph���xu%V���]� ��@��cV��=?� g��\�"\4�|����[p�e�B�{���=��f4��������TЃ�p�+(��;�l���
�$�
�\.Q@����V��3/"��i
�g������1��s+e[�;���������{��@����B�u��{6:�R���@*\��炄#D�4��2�M��<��t>K�5M�����z�t:HR��i��pG�U��_����j���۬�4%2���*���hY�>z4�[u߼�r�M���p_���?ؽa]S�6��I.�ڌ�
����ۚ��~�D:-��/�`�>�͔y��7�3wG���������&5.���F~��.릙�O�A:�r����,r�R�i��	h��0�1�L�O�ޕk\rn?���/A#96��F������n��vv9��I��d��p&9=�*w�q1$������wǢny_�[rQ+���!�N�y��Z��v�_��&ݢ�!�?[�8��,�#��$�ޙ�ύ�t��f��S���ˣخ_�H�p��@�XE�ֆ��T�?�����c�wM�s�N�X�x)ľ�!g�7�s��(�lO�0f��u*��x��*ux�u^��.a���k���3��JQ�(��
H�V��Zf�I�������R_;߄�&�Z��B"Uq��i4,��g����
� �)�Y/���bK(ʃ�E