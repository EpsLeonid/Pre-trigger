XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.*�����4e�8R�x��2ƫ��"|���I���82��$1O���E�LG8y 7��)���i�%{���̪�^9�3���Ȝ6��/:y2��&׺i�]̏�p�G�1'�>2	x~�̴V{��8G3�f���nقΤ�O����*o7�����	ñz�cJ�ε��r�OlRsD�^�3��n: -r�=�Oj���ە0��Tu���d��+>jw���e����6�f��U��$�ie�����];����ʒyHDK�i\�>w%��9�	&8�;b��-́ZU^ ��P�{�H/�b�0�a�3���уb��c�#/6������/n�x�,Q�������E\}��0�'�:��K�Q�n�S�>l���i_.�)���ޓ]�H)���'Tb�"�,�l���S4I���R���6�ϘIO��f�z���a����e��K��籔_勵�Z�%�'<�(:Q t��g	�L4�61��]�ac?���hc����@3��;��,�ŧ1��~ĸvW���P*��yC�K�G{��cauFh�Z�n�4Pi��������귂"U���q(C�e�B��@��qa���{ER��r�`��i�*���mC��!�v�amN�Ds7���	,��o�����{�.��?GA$d��[^zѴ�;���-؀Ch8$�nؖ� 'g|x	@V�3?'���E�� ϴ��R;�T1����eU�W�S3��s�_<�_VS��ts����Q�,��O�`�XlxVHYEB    19c6     900�&��5�~c�� :��'6��e�4U[��#�<�y�Ș��O�m�EUx%��][���rW}Dl����GzLaۤ�wn�%���z^o����>�`A�c�5�2�μC��9
�a^����5�J������0C`-4�*x��M|uvй��v��s����f_ĵ�!��F�1�x%�Y����.���33�.٘㑯ch��<�v�>a�G=��ݚ3��D!��&ץ�5A#-�J��u�)~��[��GP���s2-;�0=1��w��맾�(.�E��F�f$R��>=`Q�%��t��|�^;Y��7�1��e�\�c]jB�<�]��ѝA��S�9�q�P�}�v�Cf�{M§競R/��)D���	,ISՋ�^]p���^{�f�yͤ�����+`$7��\S�����<7���Ƿ�!o�!`�%4�?y$�V	�T��m������a�\��kI"�=��_�>� 9&�[[�՟��Y9Qz�b���ɳ5[�C=�+�!��1,��jGUh9ϧ���M(,h�!�h��/�� �Wi���gDy�Ӿ�������J�l]���Yn;���fһ�o�S�����R%}�z�~c�U�K��f�xj�o��ٳ7B�Igۤ�G����T?������gǻ׿i���*�=FE���6�p���;/`e�b��n}���2GN����������i⊞\��y˫W�9G��k�+qVEC\���H�	YZ�K�Z�3��n"���V��x��M���cs1Gk�gڋ�hr(|Ὢ:�51r�;�b&�G��.�KY8-ס�����j�7FU%�,�W�;�����v(ª6����R�QL`�I{�@����=ȀHz��֐����7���TD�0�w`N���� 5���4؇M�aM����=X�ed�k�j�-H���,m4.��/�ᜤ�$���y�▍�ͫ�M�?��q�w�������^����[�~��N��1�����q�V񷬱�|&B�Y�������x0:{���	�W+v������aY�H	!�K5$G qL7�r��l%\G�C��_h�!��0������p!{�)�eB��@�g,�ٔXKlV8�Vxn=��)4\ѩ)7=�ڤ�"}�x�5����4�js�A#\u3v]F�"��9�Cr.�Hg��|5:s�S�N\�+2�R�Y�s���6���(j�@ ��`�o��aC@:?U/筐䑗��+P$�B8K²�"+���g{*�`�=Ȳ$2{�7��m=�̾�>u+2v��,��&1�Fj# ������x�`)��݌��+�X�������o~��*�I���uE�VV}�7��;Z�=;��Y���vz�Y�Z���6Eg`Zے��s�I%�NQ;��Ά��?�nA���d:$�d��lt1�|�K�Y�̫� 1�����-�J@�V�լD��ThCi�0jk��x3��H+��d�/���ݫ鑪[�{��p���a�ϵ�'����X�e6e)�A��TK�bw'%&����X^g�N�J2`���(*�pHjƣ'~	A�B���`����\�*�s	�f���&reħ�Rk�֧/�2��A:�X��'{���&������y8|�$?S}�^J#R��9T���n����m�^�q,�1�U�6�@��q:���{UM�0� x[vA����aD�3��Є�l�Ì��бuuǥ��L+%V�e�u�k7E댗U6b+�ߘzQ�S-�4*xF�]����#�3vJB�:e�g��h�� ���i���Z����哒 ��K�(���Y.:�UoYVK�_��C+8��}g粅�ߌS6uz;g�F+VQ��c�4�����zFSߺ=XizZ��O�"����qSj�A9�]^=o7hJ�Y� |���L�i]^_ޘ�T���6|F��沒Z��a� |K�]`ܚ>C�U����	ѵ���z�ZN/<A��$>F��X_F���B^�.��_�+�9dV&�?qUj�~�ðU"'K�P��}RZ~�)��2����:�z"�)i$�j٘&�����c*������oA-�>	��n�#�Ц�V�8�r����3:� �3�^ k�ccq�J*n�ꇂ����[�0!���%�t��\�����?�Fub�ϞZ'�z���*g���{^�2أ�-Ũs��f�	��32�X*�pPP�.����ve-�
���Ĉ6D�[
��1��A�wZ���������Z��il9y^'G ��:�=!�*��^�������:#����	:g�|�!