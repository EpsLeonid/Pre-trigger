XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[C٩����7Ć����j������ ���%%d�p>�Oia����#by��ܽ.�W!�c/�G�S�����UO�T��$�w|��ǅ36Yq~�@����~�	<34&�aq^�>J�'X��Y<4�'
��V�h;�rݩ"P1�K�!�_US��Ьc�'y���ѽY6w��n&r�xɲ1C������1y�b��^�LHh��6���ȓ)����^e����b�Ys	�4R5������D�Z4�t�T����>8�uՆ$n�a "�<�<�Zp�_
[�����]�����~I��J��~�l�*22��Z3<\`. ���5TT$����*f ��sJΉ�"
��{R-X��k��&�۪�������懑8N��z���e��8���W�������p0T�D76�k�5�Q��!~���8�%���n�|�b��3El�<�DJ~m����o�L�~�I�hXU|ɀ}�X'��ɖ���b�-=ch�X�"3�t9�6�*�l�8u
%Aۜ���������~)֫mo%M�>���g𑓹�\�.��h�0:�9���5N�s��1a}8�)��%#.R��Ģ�_8x��w�S�Ix��&����������/	Q�PL,�0�T=�"��~�r�������l���/M�z�0��6��2�o9�_+��}c����,(_ y?v�L�_��
�|R���o�$I�YMg��c�X�߮ ~�5��)����_�gM)S!͚�������i� I>\[?"��XlxVHYEB    203f     a60BM�b��a\���|���������v4(��x�7KT	����)�'�xB�����EhÕf�_:x��>X�f��f����ď\�O�AjёЖ��?+:�dp�=���̓A������
�{�bėz0x�Χ��ǎ�T���	܋��$�_X�>�ٲ����	�Ff@ݟu7�s�1ϝsp�Z~t���[)9���"�o�R҄�J���c9���'�JuX��3��p�G[mRGc���=u��g����b{�,Ou�2��1u��Cr�>��,����M�Z�mw&~f`=@�������#��b���(���f��V��`��	o�Gz_�f+B���~qpDDE��E�A��uo�����{���J����?��%���4�oz�u�:~��H�#���/���k��C��Ko�v U��D�������U�)�8�P`�ڲ�ЯX�_A�Rt�����o܀k�N`M�V¶�)��79vQrfj\��r�oo�Կ�$͒��<ҷt�(>�9����vR q�^�a�(lXj�&�(�Z�u������?^�^����Ծ�'�倍�S��� \D:{�Wn�y��O�IH��b����7<,��0o�e!6uϏݎ��8���L�GP�|�@~v���βu�v���~P{#ȡ����,*����*3����S���T�� z.7C��������#"�'L�$�R���D����A�i�i�N����^�N��f�����n���޳�� ;_�Q1������:6D��C`E���>���b�1�{	�++��C\��~j��wW�Z�X��t6������uY	iC�d������*�MWq*�����)�����|Nz5Rq��Ǟ�x����jDάG��p�Z���e+���k�a�:����y�Q� ;��+JCY8[��O��VL���/m� j���/}`rb>Y[J �+��QZ��}ةnFM3��M�*��y��&s�9�OC����YL���өA9�4'�� ������C�{�c�����'�&W�;zZ�bz�&}r��`*_+|���D���>��7�AI0$��U�M��/v�JNGͼ�-ƯW���2��=5�}�:����*�'��� xikVy�5� 6���6�g�G��*{�v�A�K�a��e�;˱�;8���#-�^�A�v9��L����}V8N�Y����CK2Y^�|���ɩ�:t�ru1��f(�$�d�ۜR��Z���l3�)�	_��uˌ�M��Z���%�>��5� ^��.r']�k�� �)�%���'�z��<�=���q��OQ���+�Zל/����;�f��h?��a���ހ�O}n؞��Q�	5�&�Z;9�"T���?���ǚ�p�OP?�����k��i�n	�+�N�������y^Db�������w3�J��(��I��V<��ӄ��9$1��^R�6z�ٸ k��lQ�щ��ݴģ?��jN�f�٘���4�%^��`���X�~�6�ˣȿn �b�u�q�y�yC����b!�)>��yr����Q
~#\I^3pwmr�@'�|f[�����yz�d�����Ψ^u^�/#y4��J�=OГ'��~<��2��|7;�m^z\G-ɝE��`���*Ōa�\G�+�a~y�#�4{dTw��/>��%�Gd$��9z-$�G^Elb��@���_���-H�_��������һ�`�i��j��o-ft���]�+�ғ:ʔ��#Vշ��<�oX�3�x�W��1uP ��@��4j'��Pf��^���e;��$A�?�Ԅ6 @m�ue;��MF}A�c�(A��b��rrU)�������sH�֚9�6w��k���,���nߝwc���]�<�5�V�>X�-Lc\���g��/pu}ojD|n�\wm{����v�wܱ
`����lI,Ԗ4v�ѝ��y{&�xh8���djla�eG��-8e��H��1L�1bʼ��8#��0�_+�H$ȟ�^�t�xGQ��������H[s�y0�=��$��@,a�oq�ɒ�]��L��nd�y��A�Vy�i�2�r�>���T;*!}
	Q^}ԯJǥAI�E�����'�e(XW<]�ڜc���,ɓ	nآ��'9$v�P�����u�� P����Y�۴�`���ۮ�za%��R���o�����/�A��{�v���:Y�/�Đ����j��ּ�g8���ŵ��c�B�����V�<��*�}/��U�im����������ẓ��WW��?�����+��!��@��+���ki�(�-ΤE`V�<5���@τ�z-�6�N�|�l�e�0yD��ٕj$!ChV����V2�4$��OP�%����L�)���aVq��#����&ܧU��J�S�����ܹq��6�cY��y��ZR��!��mX�!�q���G��T7��[ �Qw��p�?)u�Q��Ld��3��v��lCz�qЙseH�:��!H(�=�+��U�-�H'�,�B�d��=��B��`��N��i���W�U$	-{���~u�"M��c[����4����qs�P�lCm'yA"\���G�`^�f$7�.�GӘk�:V�2��9z�Y���,��� ��Եh�0��