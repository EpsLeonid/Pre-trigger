XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����̗���}P=Q�g�ۼ�Ȝt�f�8b����*g�ʦ�h���rGA;��N9>{��^p�T|�zr�f�v=)�3�6���1g*��,��"߉�1>�P\y{L�0ɦ��i��7B�Q|��@��K�1M�dP��u'��^�#gY�[I�����@��&�׳yf*�s�*�5�<'w�#SE��@C�v�^�(�,m�v���A�L>��;�����~��#��ˎ�D���^�n
�B~XfJXX��i"tC}������vߢ�D�ŗ�Dz����YK~A\+��j4�z��j��i�U�����P��O���B�c�O���b�9���!�-R�9�>�q���3�;*"l<XH{�� �"|��l�?��"�+�w�x�jɢ�i�ѶW�U��^L�u��@��b��gD�"p�k�S^Z�شfA��(��Q�<��%����]X�K�X�A2�0�giE[Q�r���
9���2�8!?�=�n�@k��B�n����W�LQ�y��%��^f�i�y\7>��B����Y�-Dk��71�C��,�K��,��p8(H��=pȞO��[��J��":������#�]@S�EIt��I��*A��R�@�ݒFM0|�e����f�)zfϣ~Da�$h����<��j�n`�%C����ò�p�:햞��Us�g6�)���I�����a���\���#�^A�;Mś,���JK�u'���<�LY�����֎�� �� �|"���U��] ���|):�_XlxVHYEB    118c     6d0�2���Gn�[�M/��3|�y`X�%�������c�ȇ6�4B�!��Ɓ���d��؝	.�j"�ā,a�4�Rk��u��X:d/1ȋD�WT���/v=+٠���*HpF��֠�P�+�����K�uB6}���{���Έz%v-N#K�o/v�;Zu:�*?Q�~T�kV�H5a��^�4B)���#2��(;��2�J���|�1~
��%��c���I�֪�a$���%�a���oS�EW*��/�;$���u<&d�$����B�8;��h�m��"�^�ᗆ�"9���N�c��j��pXA�	���2+NU���[��p)r�.C��Ϧ8+��1����م�-S0@2�޲O-�&x"��]Pdv�2����?:�`?�1e��׷diq�^��n�}���
X��8�ݽ� Dw��NM�0��sP �K�������?	q��ǏGL,��	�J���M��z�I����3A����t@�\�����A��4���.�a/�M>|��Sr��:��r���rM�?贻Y��,�����Δ U�Դ5���;��=48�l�J|k)+�]c8
�QfZ�i*r��������?�,�����':�>rǳ��҃�H��<�/�eO��Z��d��A�B��t�ȯ��X<����zQR���ض&�_�U���-(]I�,��<�j#U3����6+`��������.�v�O�M���,��lO�Z@B˚ic�Oy���N������G���WR;vI9��>u~g>(咘���t{]G3��n��t]R��v�Fv���+�7�Io�����r��-?Y�Z.N<���%R�7�3i�ƐT��(jeo;��Ѥ�l�7��.J�N�O���A
�g���*����(�D���s�cs�=��/�G1c)����q��ϫ�'�����G���G{Ɇ�GK�6�xteJ_Z-: ��s;��Nl��71��Lʥ\����҅�� �9�?�nIj����)s��D���mf�1;�����ӳ��' �g�eM.���5Yӳ@~SFs
<����;]��Ro^�J-Zg�}�l"*�F�c�Z���?�?���1!�Ձ�eO�ӡd @j�V����	�fe��.�xv�%�&6��
�8B;��P)�ڠ�����vI�����E��(��c+�>��C�
��^u������G>[�=�Ban�ů����
�K!�v<2	bI�-��omp�BN|魫�Gd.bc�OV߰D)�3���js���F��XG��r���X8�F"�-nM �t����K%��{b�0�@ås)(����A����e��o᫆}7iv2����]�*�Ǐ	)����<N!D(=ء���{���G�ȏ�X���T���<�8�3w_�1��+�t��F��%����-��q��	��T�����93K�+��S��U(�э���x+P�2�j%9�3}}�cR�lM�I2��z��s��C���6�u D0��˳��!��@i����_�:<�e�|����A���]�x(W�'�[��~R�PU��N����,rN�޳�
W�S)N7�n?��7��	[�¦.)����'��(�Ԍ�/�2�Y�\e�Mm��-Z��?'������w.��a��|8
j$YV���ϸc,w鴾(����ۭ��6/��?V�N����Z/G����7�