XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��؆���h��Oꉽ���
���ޱ'P�{ye �B�����щ�x��'R�Z�r�0껨|�R��#�Rw���op�kһטؙ��߇rިP�|���p��߹#�p቞{u����e��`���#Q�Ϲ�8qe
�F����8�B[���Z�cu�| �����N������UJ;�|��/I�_'�N�'�k�e���S�`�Yǅl?ő3�W������S�8٩hb\n��b{Q�X��6,Ys���hg8�ջ4?�w�/�U_� q�?�P����8���)}c1%J�a��W�)��#�
S8���г�(�t��c�f�0 ��m�7��f���)>ׄ���c�ݮ#�O���6����ZE��,��*^�c��Ǫs��s�y�����>%b�
����I�d�C&��S_R��V�_���T
�_v��1�mwl��]�J�І��c���J~��pm��gH	�T]�(�Y�����%x���v�%0{D��*�������T;%�iaQ��ޒ�q<�FWu�z�3�/U����^�t��
Sl�n/]~<�d�Z���<�Pr��<K���m�s���J��x�G��2�Dg�;t��U3���ō�y����A�xMgɼ��k_�
��ب��G����p�k�Q�G9�0�6��*]e�A�]���V���)(��5�5X�����*R���q��bq+�e��W���_�5�"�U�x6'��j4�*������%�5�{v���+n^XlxVHYEB    19c6     900 ��s4�I�l�fKN�3��
32H�%X}�b����7���g�v��0TîJ�0�3$�rk4�Լ� w�G��?�\���D��i���N���>����L�i��h9ʎ ؔ5;����ƨ�԰�ETpo�k�����y��y���ū5-~k�g��S	z�_;� Zo'�_>�r�И���O<1�V(�w��;��@�ƢP�SRjb��'�X������h�Gz�|vu<V�W)9�\q܂W�G���J?�GP�� }��hQ�N�"���V��J�����Ks�(��Ʋ{��������S�Gx��C��I l���8I��kh��.��<���`=&��-p�ݻEԢ&�ϳ&a��qE�z���d��NE��Wڐ�Z�ϼ.<�2#�z��}���9S�y�����j�sՒD�/$\'s�ؑ�ZYv���-$�q@0�%""f}�$E=-r�*j~L�?����8�i�P�n�*h�b[o�]���l�~���\��mbw�ʊ��[�i;�l�g���qDP�լ��,�MPo�Ė[�ް���F�3�z���&�@�s���>7p= H�q�죆��PA�[B�J��8���t����WZ�<Ȣ��y럳CǫRKʴ�p�w�qn���-Zh}�-d?��Vy�86Ū�XW�5����}ᐃmo�+\��Ԝ�;�Z!P���t��!�qEu���F�����Z1��&{m���/x;�c��`��ڊ!���<��ӭ]�m�u�dLE��N��& �6iq�K�_��=�d�:"1:�M�A	;�[�Q�4vQ��ɢ<<p �{�[�,s����qJ��S@8�=�xu�k=4�EwI�m�=��J9��P�w�5����r�+�6$8�[��h��$t.�a�������Zɞ3_\X�!�?;��3c3���Ā4G��<��jO�	9b�(��� HS�Jt�����&�Q�!��1{梕+�lL��@�G���X,bn�7�r�7<4WX�3�+l3v���Ɂ���Liz=)���܁�dq5�ɾ��Rg�9;���n�E�I����dw�������g7y$:I��3a,��{�a= ��_'��0+|�j�/|��	��ŉi'���A'�&��ˑ�#p�6��L6�62j	�nO��o�."�oz9-�&k�j��)�ή��+�1�^k%��Nhis�:B|g*+.��yE-W1��zW��+(�q�;��J���5˔��H^���f�A�[�-�!ߠ�O��w��n���*��y�9?7{g����dr�Bkʪx-���B��į����M����?3s[Y�Ts�`Jbo+�̄-*qXBE-D��μ��Ѥ?�N;���i�F�h^�,|�x��0d�S=��.Z8W�[���_-2z���s���"q�V�md���',�F��K��G>'��'�}trB`��j;\���(e���1�a#j�~�2���t� [}��g�����Ս��2>4�m�7��v�V,4���.�]�Br# ��j�K�4U}a�V���zx�l�����`��.86�PB'arK��[h7ip[Ӭ*9t`u��T����3���5��6	�f�x�N����	M���ĆPS� ����g^�d��'=~��!���@}g����mK��j��ha�RH���g]qp{�Ea�����~#��Y�2>���ଛ�*�&fɧ���>��#��H_��$vY��i4�7�Y�( �6ΎY�g�H^�"μ��q`��/����]����ˋ�ې8v5^�븹�k�Z��޺�m鮨��%z�b?���N���X�@�$��+|Q{(��4��2���:��ٽ
Kt1��z6h��D��`	��p�F��KPB��	��SxXg�ZG5�N-0���o���.8�%����xv�*w���$�8��e��0o�Iq��՚\M���	ϤҒSλ�K�	7BtK�b�Z�S�5z&hE�x}[��zl1��\�2�|:0<���C���wGS�Vom{!��ټ��u.Y"Ό�^���Ov�k��J���?V�{V��߻�9�*c�3+6c���K��/c)ـ�q��	l�Ga%#��y$s��;ĳ��C�y�Z�h�^���#W��:e���Ş��[^�ߵx1^oS��_)�Ŀ(.n��BG����
�G�{��=!׭���?+�Wp�	�o���Y\C`p�N��)D2�E�D�~p�ǝ�I���^5��b�b���/�\e ���v��q�yo��`�Z��4'd��&A�LWu�Z�~&�-�gv�T�«��