XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P�:��d&.�f*<}��x�� 6�0�����U^��E7DУ;��!9~�vV�LIpV�+}f���������� ��
y���v�7⋚<7x���\�>��>��}	|�j�K�j\�EZn�b��yXF�;��C�����T��J��B�9d�MkP��t����Ue�_Ӊ8�".H��6�����VH�6�SIQ�C��k$Ȭ,��#N����OC6�ݼ�Z��SO�JQQ�G����D��GS�ͣ��p�77x��V��B���G��^����k�:
�}�G1�0@���I.��)����\&K�기����wa�¸\�ӄ�����u�g�����r�Ж�����sE�%>���A0A�@ O���� ��QS�`��~^�B��2��'U�v�0�AI���~]����(������d�D�wuRᩘ� r�v �$��W"dr�#���cCC��5Iq�o
�
 �}\y_��[�S�e�F�4A��ev��J-x.Әu��LD��t�s��I�*�}�*�K��J�������7��M�!����s|�&3{�_K9�ԗ�+�Vm���7��u��]�my�P��6Bι-�cǊ��n��ɡ!6�
�� 8�̋�����g������?)t\��"&�}���*D 5���,�s_ܗ�4�M�b����˺��Gc
\?
r�t�����Z<ﺲ�����=��9�l9o��%��2�7����ܗ�,�s���_��UY����FKXlxVHYEB    1a2b     8f0?�hM6_A�2�k��~dZ�������o��=h`R(7b(�l�#�����%�X�9i�[a�Q�W��.A{�s�75�<	�
>dK��0M���'�FL����u5��Cm����$����J�n��Ɵ�;rz��zte�Q�>6�^��S��7�tV�mY��N��=��xb/*�\)g�e��~~��EZ/��]o�b�0s�P�^�� �����C�bǞ�-���?�s�!ϙ@u ǐΎ{񂌟��[RW�=��4:f�[+#�멞��Χ�g�˗(�b�|c"��!��?��t�tр�Mo*��+�X��<�4�,g�����y�@H*^���ͼf%��מ�W}诖B�ּ��N?*t�}8�6����>wY[@����*F��(x:�i��(�>(>;0��!�ES�����o45B�U��:`�&��;��6���&�_�!
Mm	~t�=M,_v�+N�� �e���(�ٜ�Z�X��l�7ϘF��S����糁`��?o9���u+[^��o��I�n G�GY�n ��sK���X#���ߪ[�tn��ʱ��S}p=|��NM2���C7����W�y&9b��璉�c�LE9� y�y=�hi�YH�~���_��q'��m*Ο�b���H%��M�u�&�i�EH�Z�밸�����zHT�@	�����6��%Y���+W�t���ۜs�3���kUV�D �	�$I'Hŕ�������K
��[�������#����xܼ��7�K�d��$�\�!j-�+�ע�Vφ��>��g9+CY��`�K)`�ݟ�nCH5YT8�a��Y�8T�2�9���Q
��x]ܯ��/]݁�r���¶�q,*�Z��a��޽�(�ܻ�.��'���?�ʰ8L}�I�˜��R�kѿ~�f)VD&\�'Б��40�.���gu��Y�}G�e���(g��F��b�>ud�Ȭ�׃���|���7�W��j	���}��g��62ىK^L�����ؓ,z���ÜԢ57 `���T�c�`s#��?؋��:.�<)��{��(�$D3ᇮHx�����_RZU�S%�i�}q]�F���,�/i�>o<�Σ�K��pZ�K@C@hdι��,S<��L4��`����'(6�T,ˇ�&M�W�^�����-�������J�[��YP<H���_wH!)�p%�Rv_�le�$���::w�Z�G�戁���M��O�Zv�C��ػr/�<�b�[C�x�@���ّ�v/j�+��Y�7�����ɱ�U%,8������2�� G�J0�q��&6V���s#��y<R�s4vc��0�����!����Ӡ�S��(mPM[C���6�RP�_����s��(�2"h�9�ӝ��k�()&�v��8�R�O?�Xc��t3^]1�X.*:JU�C���=���osE��F��pӬy�N,���V��3����)�U�C��w�|,�ѥ�d���L�Y(11d�ɗ֭6&"��e�M����������>1h9�g�E4�E\�w�����@B��a��Pn�ߧ������A0g��x�KՇؘ�!��i�-��d�0�_�珎L�j�̈�Y���ÍP
Z/�Vi����ZP�"\A\G��f\J�?�K�X�hٲ�ce����c���%���c�3��~O�0ay���s��З�'�K�q}S$���tI�O ր/�,��� J�-H�y�،�,�nNl�;S�π�T���n[��M�%���&�'��r�l:�:q?}������1٪^���eS���Q,�����S����=h�l�����9#�OQܐ1�j�.��0��؁߁�'�GQN\��y��_4�M݃4��'�c��չ�UQ�b����H�U L�K�!�?�D�;�0o�˰����Ô����KmCӡQo�$"�>G��|i��&?���;����z�����X?�;8m�fG���]�D�+P��e/��{�Tt�+Q�����TJ��?����N����m��g`D�TT�[�a��7����8�YaL�?�ʱ(Lh
y����Ҋ8������oiQ�B�?�����b[ȟ8����%��v�!�/'��d�>4�}r�h:e�D����+>{y���mv���o�~��o���4'[�*���!��h�4�m���s�^��r$�ҷE�L����\� �,����ՠ��~��4�
ư
h1[c��Y��_&�i=���~��X���FG���Ç1��	�~��~��&�����E�]�0q�