XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��7BW%xܦ�!�u����7'��&�;�g�]��d$)���o
�C�k���O�^	tdQ���t_�j��I~�4��\j�9B�}�BԎ�/����g�~�F�6�bF���R�w�F��R�WF��;�p��+����i�2�IްvV�m|�&p9��9�v/)�Y�3ce����EJލ���XQ��m�s[���>�6�}�^��<��]H� ���.���kv�N��K`6b'}G�b1Z>��-��6����~��9x-&e���DS�ز��-p�#Y�G'7�)�m)�n1� ���]A�߻�kG�lRT��ӳ�%09�q����8vy����VW�S^��j�	��&rJ��L�h.�T��p�l	:I�U���S�����|����=y���
�־�y�1��>1dj�֒B�
����4����B��i�S��$�Q3.�>�n��;�m�IF{�禺�}�=* ,�?�V�P]����c�=�3g��b��v�)_<��*��`^�>��Nn���~ t�3@��]�R& }m-π��H��&��J�H�ClG���ȅ[ ��Ԅ��u
8y.~ڀ��漖��d��F� �q6a��v��4o��	�S��Tt�B�/�v��ޭ�93������~n�߶0��E*8558�A�=��te&�@�~�?�L�	X`��vL�X�tG�QT���2�ԃI���*��� [��(��׌J��L\�9�]6CM0�Hr])��������j���XlxVHYEB    3292     b80�yb�NF�2���h�2����0���c&x��.B;��+�rE����C�U�?�э�:2RҔx�����.�����ې/�4��,o���ӝ�m�s���x���]��n�#e7�A���'���sa7�I��2��Ԃ� ���;��bR���n���ڹ^6�S�׭ﮪt��S�
���b��,�P��\���<]J�Rt�4p4�=n�~�'ѽv	+�{=S��ぶ�w.m��%�ׯ��y�_��>�k�r���%bP�MW��,z���ݸq���Y�jM
�K"����w�R���*Dzt�:�����W�
f$�<��.��&:�3]-���+�36ͭQ�;�/�9�<�nnw��=�C��8���r�A��͹�;(�,6��J\��\��Uj���B�P'���eN'#ۧZ{�8�<��=藂�M:�SVwP��8o�:�����O����)}
8��SUg�=݆�L��ŅBt�=�Ӟo�s�����Ae-�@�r^|�X/����M���ʌ�o�?����U��T������Ү��j��`ެ���,c匚��=L�D5�w��q�����hu{��z~D���� A]l\�]�M-�� CK/ϰ��k��Hy���A{��,a�{K>�@Wpf �����]`Χ4�m2��Q�ݕwm�)e���@5���n假�8�mu�9^u��m������-����hl�k;��
Z3~��s�Ѩ��~�����+��l`�|�U��� �3�Cc6D"S�[�:���>V�n�2\�_O�'r���LC��PcV�ʅR�~��O�џ����2Ӥ���X&�!Q7���&�E��~���t��m\*ig�n@p��T,VPrU�*Țv�����B�	QaMj�Np�9���W�)�ͭ."#N�o���.C�+���_g����O�B�
$�@v�ٮ�J�xBU�'��>9D)nDM��|m�N�L��1�:�DWZ�+�9�"$/�>��[P�/r�2��8O/��\\6��B.Fm��%�J�t�S|�:;����U� 4ԋHZǢ� ��O�k�o��{<��>
�@&P��ꃏ8�S/�zJ��lpુ�]�z��3�e�Y��Ԏ�;����M�NaB���,���#��Z�b���#!� 2wS�i$�ű�̙L��?�qm����u�ٍǱKS�)�n-S �'��(��)���-��R�8ۘ�A�:����\Rw9��-�dX����5����/��0�D�4�p|�N�Gp'h۲x�NsfF8 �-�8 ?e��`�K��"A���X��VQA�L��������jv�ex��IN��:�Xҁ�4UZ˄��ě����	H���2��Z���Q��$a뷏0q��U#lq����]$�(���Kk6p���B��+~��	�P�'.L�F�|z.,)�@��?/����V���_��K��\ã���@>�}v���*��YgI�Ώ�)7�a^b�Z0��`>+ߥ��xp��>f#����VO@���ɔ����FD�<G,3�;䱗�j%�`{�9��	Ǧ#�W��'O�]��%��񎑂	JR=�P��a�ʀ�Pɍ�H�����M�W#�u6h[��GvMg̠��r�5��Ep,WYX|����#R�X�����;S��}l2�P�Z��~6_�B�(а0��I	&�h7��\Y=�`/��m�>���R���Y��P}C�ǻ�z1]���]�]1�x�;3
͡`�� �9�w���5nAQ4@7����.�m�F=�*�Z�F�v�7� ��$������K_��зv����M���\�:a&q��N"���%K�ˠP�̣]��G��f�I]^�i��<�㡈�3�Ր�KK���V�2��?:S��D��|�C��mFp!�����܅*�x��y\q�������k�y�� c���1�Uy�m��v	X�����`Q,Ve"k<~!�|�(�FBrΈ ���K���A,-�9��	�u�� ���j0�@3��y_Jܧ�����Z<2[FL#2b�
x�&Z�d�ɭD��";O��3�H�
W�:�ݞ�@qȜ�}�1U'}ǘK[>%�^���QXr+�Ȑ��N�F��y+G,�w,JW���{�M���H�d5x����E�������Yk�*�*�+��GQe�O/����t3l�,mp5"�@��:[�
FMiyɕI%g���h�"�Tp�
�` �֣5K%hC	�!w`�S B�с*�*���b��������;��I���b�!��?�MF1�$D�,��)�ݼN��C5X]�����;SB�MMm���:#�f�]9��GL�� ��͞�l�/A
��D��A��@����#wwg�x�j�XM]���,;7�E^8?sX.�����֫D=�I�`\�l�@p�Ƚ)=K3ùʋ5W��A~ґhi��[@��ch�TU�2��|��g�.2M�H�g�:����U�P#<d��
OS��Ϛ��op���	ﴒ}M����)[+�T ��\:���]�i���Z��Wa�ԛ�Z)m�)�QH����x�߬t�L�
<�@����J�GG�� 0���$�ۖ�2���(=�#�����h�U��u�{y���bF�2�'��@�U䍤�u�I�V)]Ŵ��yb���gv��bƦ�����[IPlm#b��i��s<��}�Y����X������**w��/\��.|O=��"W	�V�0ks�=�6���l��%1f��<Z&$\�0�8�r��G�Z9J\kr7Y�>}�������ǲ�vd�݃�;åm�� HFG�m�M
�@�� H�c,���0f����r�om�qޯ��������<U�0$>��O;���JF���9[1�I�M
؜�\������k)B��0+wZ�����~�Xh{ ��<'�Yqa���+aQꥅ�˹ۭ�V@W�*$�7�/��y��u[0