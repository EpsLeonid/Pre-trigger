XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����������������$�^ϟ��/�ՙ_Vʫ�l-Us�xM��\���Ǧ e�yI*`^-_��=��[������(2�L`"�h�!�J[?��b��P �G��(�q��#��AP�u"&�..Z��xw�M�6:������5B�� c�������ۺ\�}ц��0h��p�P�f��tĲ^��� �T�rd{���_�
�Eu�A�MP�dʮ�P��+g��J�4�1A�^k�ˁ͍4WT�e�~Y�x>(Uތ\�̛�9������ύ�3/�RQ�BwH:	������Z��s'�;��e&�W��:|���t�C:��8Sg	�%sS����>P7٬�ǚ��ه�F+�"����+|�	U���c�:�`���j7tz0��
J�E��(k7��5s�K�zM�`a�������Ȗ^0�$���t�����V������K !�
M�5N��.�e>�#���$�M��9�o¿*�i�'h$G���q���8��b�Ot�s}6B����>ϰ���<�������L���D� �*��C�l3סfX�I`��ƾʧ���[����@3��I�8o��+�%*9v�*�#C 	X�|2.�v%�]v#C�)p�5�ZX���e{(<[�^c8@`��=|q�>M��S���:��Q_���ubx2�Hj{+<߅��YCnk�b��%��B�`.z����B!ۓS\�Z���<�����گM��V\���g�'qU2�dX��uΕ&D�մ��k����DXlxVHYEB    bc57    27e0���Z�%H��3	�j1�&v�?���O�8`�,��B��-<�����˥$EªZ_�-�b�>	Y��	h�c�gf_��J�1G�Ë��^��Y~Yv`�)6��ZYp�=� �����;�+V]H�;�F�3�ʴÆ�:@�bP���Ʋ|k̨����8�:�ZT?�-��N����b擂���e���}M��UC[���%����'Tn%N;�9�:�zʍ���!՟r�lr}��G��Q7��]���`�l@�Qi#�
��?�o��'�v�}����4_��/=�y�&d�1dAxP�7xx��1pK ��F�����	��#����-e��qB��n��/_�����Q�ׅ?
�����"{;)#t�ay�%�?�ڿ�56 ���pӝ��"�����m+�u0B�H�yjL�		�$�tngֻkh��u��2&T=(���f��g+������z&�>݅,p�<�(M��Ⅷ���3��ag�
�2����ς��Hf�_�=�T6�s�)�q��-T�k�rj2Ķ}6HH�ŏ���a��ʖi�}��f�݌����]w@������A�`z3�(^����H��I��	"P�j䱴Ó'���[ΦɃ�c��R���F�_��C������9��,vh�D�������0��I�q�V����S���It��"�u �8D�v�>�ܽ�=���Y�D�*�vAQ�?�������N67�>gP�t�3$�]�&��������p�>�V{�������&B��%�BA��8Ha�F;Zc�]�x�"X{��x-�7�Q?A�����>�9�^A��5���;+6�S��|���3(�B&J(���=C14��U�o�2j�B��[HPs����P̘�ݚ���ca�y�zV����x�9.<"�������*������,"�3�ݤ���qJ��s�UP�PK&��:�f\"�څc����N� ��s�JO�N��w)$������Z�ϼlY�����Ai`��_���S�(&5�M)�����?"�^�bx�{j���t^=(N��8��j6�����2\=��Cc����		�:�R���� ���J�bķ(N�e�D&;4�����pՑ(#��;��P���#��\e��u@rt[&�;Jj�[u����ӕi����Bv ���]o���%�ZF�Sш��Ͳ���~w���ǳ�E؊d;m��*p��(l{�Z��BꜰuR��)���}��^V�`��b:�c`x��o�爷�Zp�%w�M��9Q${
��q!ù�Co�N��}��!y3��
�|/���V�^���
�"![���m�A'�FG{im��8���_�˴�+m���D�$����Č�}�#g�y�,N��,Q��,Qv�f����]�(?e��sC`V�:���J6��R杴����]L$�Ҵ��i��L3�ǚt 4A΄x�8>��X��G�>�u���}ݚ��?'�H�'�un���k�ڔjă�7���%�ѕ���^��l�t�GA(�A`�)���F9��t������2 I~����"�����,1j�jrx���X&�Э�|�ku�0��B6�g>܎��1jd.�N�5�t�rQCF�Q|̎N�]��V�\Q`_hY���D�C�@kD�q�A��ԈۯHv�x�w��Je�h��U�?}T;�O�{��g�8��w�z�r�(�������#�]��5�⫥�z\Sb�/t���<�pՇ0 j�Uu��&��_���U��@���c�#�+���q�۳���;��"�w�2�Q��Ɂ&Y�&���
��'�s4V��MoE�\PA3}Y�1D�2��	[��,B�Ô�O�^�Հ��x�?����(��_��ɵo�;Pς��<��v �t�(o��X4��p�m{��3ęd���`ϕ�Ph���Lp���wS[�3r�̼'>���ŭ��#����b����(c	 ���G;�G��/�o�q����ܸ�6հ�����ߥW����^�@d�q�e��N19�s�u��mc@���?���1���Y@�wի	����:�B�oj�=��=D�ġ0�^-3~s���Ճ����18MbR#G���bط@4��s�Znfu8���\�)���4�Ĝ��9Xǳ�r�s��Lp������׸:7(=�<y�F�X���)�f%�x"�L�)W\�'��ݫ�H u�ők�U�D~��|��U��F���ݮ!K3"�I��9K���!�/
�7��˔�E���t^&[/�	(���\���6��d��V�;Y����uz�]q���6n���Ͷ=��d��+�ZVG.�Ǯ����"�ig�k�t[lZu8P��'�����;��F
�N6���	�l%�<�i��~4��4��C����si��ŀn��;n�a?�+O�j��hh&��Yv�2qסi�ˠ�vȤ�4�-�Y7ޝ९�Y���C���?�a�z)�a�p6i�Ԝ��*j��Mw����\��.G1�h�!����h�R��@����U�#"�"����LN>)�`,@`3��}�����x����e;ɖ>��!a?Ҹ��Y�ۇ��\ ��ɱ7�����3f�tm �����O�)g�D��ӏƭ��zd��Q!BQ�Һ�� !ȁ��8}�{��ӥPY�drP�q���J�;6���)^�u'%��v�E�{|5ج�_#T�Dm�}���9V���	��祔kIZl��d����ˋ��f�ř+��U7�LƩG%]q���m8�@�|���G�×�L1ߵ곥�u���C���gᨆ�l����ڞ��$n��r����oՏ�����H4[������ez���d��M��R��C���i�A������,�Z9q:tw<�0CO���]���ϳ�5հ仫]���wZ�ʖS�`�9��0k�c� ��XQA���d�n�����Z֎����H�;�JdB�V��SA�Q����Ơ����z�no��)�"���
�������ka�?�����YH-�0�p�K���(�C�k�%�xͭ|��E�5��HQ�� �A��V��&�{8��F��I�w���z���X��I��!��H��L?ȥ�]Ɓ��/����[*�Mص�_��'t��^�Z�U&$��&s��NB�����Fr� ��F�wLkeH4��������nsw9)�^�f��o���$#���:�r�� �[�5?��2>�ԋA�&��K&j�j�����u�U{)����^����XXZ
7�t�*���tBcם,��o�R�S�g�bz�(���#>���,+Ppoa�C�Ns7����X�	��K�`;B���|����n}p���>R(��<|0��c>d,V�0JO;�����d��VA�5܉�C�Գ��/`%�g�O�9i�'r_��� �Y�~�J�P����?���/lb�1nY��pr��T��W c�*�'	��5|B�!z�,{��h�����<�����=*�n|ے����zMJq���tQ|T��Cf�|�82>�1������ЈOZ2��.TN��N��[s;�mr�O�� �v�9���� ���gvʐׂ}�����|��I4���{̪�-��,����?�x7�T���_��0�ȇ�{�p��"l�e�(����/�Оs�WCo��):��4�����>��v���=n�������p.^�~��q�~5*,�!�K�,���n�;���#�)?4%5NAkۡ�-�l��6�o+-�ꮵ$��b�lEi/����(����`k�2i2�zDOAB5��}�2.,vp-R*�o���Z����M�@RVkF	�{(��~SS`��f7H>�6���}H�G�����M�bf�Fs�cYM�H�k��c���-�<!At��K�Q�|J����π����w��d���O��g��`��=s��W�&�
݁5}��CO��������`NN�B��}��e}j���H�2�c{�u�of���a�[y���
z��LN�w%���ª(/	���!2���7�������B���q�E�N!�����;-��C+��!kd�D������l�Ps~cB����0�WD�.@�8%(W�<��o�:�RH��ZrKOu C�J�=��0��]�Ce��4Kg�<H"j���dUIy�L���t���-�� ���@6�@�H!=�(;7Z��1�{�i�c�yB)�LHʽ�<��Q�NEYug�Fn�L~�Zkz�A��P��/ߗa4�L�!���i
�	�����#�3�2����4L��ܣW�~�5�ҕ�L0GZ_�C�hV����N�u�&� 5i}� [��'cI�V��{�7Ec�i0�8���&�{H�n7p��>�bMc�"P��n�x�9���o�$��A���X"r=_9L"
s޴<� ���6ѯ'rp���<��r�`�����Y��?. s��!�De���\K��ǝ�<&��p�gN�7�lv��A&Ō��	{�&�?��<�컀l���OC}n҂�OH&<���B�RՍi��1�dko�?V�Mȳ!^A�p�Ա4{,b��j-��!k�=v����O�F-t�R����M��~����i����C�[� 0�����᩽U�����!����z�~4>bTn m��@�Ϣwqf|鹵�c��FDpk�p�2�7�K�U��@:b[�z����V��T�u��h(�*DlX�I�=�)�8l���9��,��)��PsC
U	(O������������ٱM��*�b�aƶ��_��ď�W������S	�\ҩ��Ϛ	��S�W�cC��N������$&qx�e���m�ĺ��D L� ��U��Y��,4Dii�7��%���AVsG�tfۊ�Y4���p0ߞ�r����_�V�bf����.뚒"�J�q}�ۥc`N���_�0	o�ʖ�s��$U @��r�˝���-d�����UD���;{x@�w����XQj�F�y�-3I }��P�ms\�_�^�����b"� 1%�p���|P�$z�܊lf�Xʹd���+|,Ba�NF%�@'~�CH���C��4���G�
��X'�Z�'&
[%��|��>@f�J�:xQU�L��l&����	:m3�#�-�����W��Ԏ^t�۷q*Y��PD2���vm����p�c�3ŢW�`�.�C��:�[`k�)Q�w�H;f�,��]����#�YG��^r&�TV�W��8�7	d_U�>}3�0��S��e�3�k;{NE��%엀T*`A�M�4��l��J��)>��7Qm��Z��TV�8v�/>�+�ql]^�t��fϥ����d#���x��~�{�A��C˨�m�fЇ����	d4��:���b�o�)s9�	sS���(}�z�Q���Խ$˖���NC�M��|,��-2���v�˃�r��PZJ���R̆%�b���x� ��Kʛ`q���Y�i�H��T%��P �S�
��B�T@�3n�(0G���%��E�h�v��P��SD��(��3�5k�<��P���`�)��\r���5�a��F`��`+Wv)��zN�k����l�j��v+2��[������ރk�m�0�����;��R�#�����@B�3��G"&r�pdnԩ���|	����t�}V�!�Fp�)��"�
��~_���_��<� ٺ�~�ט�jk�W��!�p�m��8�W�����\"��-ͯ�:�a-0<Fo�A�M�Y�ۀ%oXz�?'H�q:����evU3�`[SP�ˮ70�@�c(h�����$���:c�������}�G�Qd��rl�L�`%�������%�����p�)���9��-"�ߜ��/TN�)�����(���o���l3A��U2��	)2:�_����"���e���R�T��hk��=�!a���. �lJ@ k�=L'�/7{�	�^���uv�nh�J�#�/�A���e0�p\z�ۥU��`}�!��da=�gk��"�����짢&<�;�����}� g^\C:�G�|(�i8 �y�����Kf�q����-?�	/�Y�J�h.��9ѡ�ڸ�̀{9'�N�qg7�z�	��!����i�ݫ�R���jٲb�Ji>�T��m�a�ig�Ɲ�Qښ=�����HNb"2�6C���j_s�E��&�f���g�v�v�OR@K�N�`h��W�^�={�8�`��>�l{>J��
�n�M�Q��H6l�i6*�Po�<?{�*ЎU������k��h	�i���j?^�.�kW|W�$�R�t�wT��͋�Y�����"��M"���ӵO�%�h���a���;�Lt�0�����(KJ&���H	<lugS�s-x��㹺o���ط���)V9�V�������ң���ˈ�Q��H���el88HG�8��>f#�����Ut%�[zdR��bmR�x��Ӽ�q�J<P7��-^���:�����>������8l:�@�n�O�������ؒ���|�Dn��`N�]�?�����*��a�-i����1���!�Mm� ��%ժQ	kթ�����TA9��`�m"H�L���®>��)X�jˆ�q"�d��c��ʩsFo�i&�lEڝ.-qtdkM��L@��UI�!߲���3$�{�Qo2����2!��OW⟦�P>�DW����F���������X[c��	����P�)臾���콾M�Z|a���"������Nƌ�z`_e9'�KP�,�,��B�:��Z�Y3�΃�E�����s� 
��f��6�U��Ɲn���.9p����+��f"���=�V}I����%�{��3(|�,���42�N��8F-	�����s�.b*���z�E&�Ղ�7rA#�ϤB���:n�����V�eM&G�Dj�~
�cw'\�����AݶI㍒����1i%eD�U�YĊ�� �������)$�1W�����ho�⻌�sֈ�E�0b4��Ho(c���D�6�,����N"�A�5DcH�-g�x��`e|�z��$ڃ��~2<��f� /?{�2g�0A ϊ��m*�p�)`코v>�&��fh׈���Y�[K.��v�شǜ�\&��n
 4�y�:�����X�i��s�H�+M��R�/�鳷���u#��:BP���������Ծ�9�6ܦ�F~�̹����pQ�oR�y�Rf�k��}ޏ�D��:=�NTZ�הJ�NJEl��0�	�Ɏ��6$�`��֞0���R��Ki*n߫�P;�2*K<�{i�2�cӠ��i)�U�$����V ɀi�ۮ���S�	l�i���`Bmn"�F�x��$����;d�\�ܽ%��gu��̱F�~�ϧ��7Yx��+ g�K�t�4��t W�
���(r��	I�F�sVW�ua�cS������B��$c�>�B��*[P����8���S
��aU��lqX��^q#۝��^Gv_"Z�m+i3���A����Ï�ڼ�q8�f����뫮�&���q�� H��I���e}M=�ǈ��]t���i���w�o���j��BSP0n܍�?#@����h�t^K7�*U~&Z;���yY�C��vM|����U�]����_Z�6ڢ:�^쭕X�=F���=ʀU�	F�[�r���3[F͡�@H���잠4�U�����̴�Il���˺��\��%��u`�׾� fyB�KJ����D�� �����%k`��|����"�9t���SX~��s���m�"��DDm�E��^���W��AH>c���{��6�78���M7�����`����F��ǰ\_�$2=r�T|
 ���l�P-�~U'��%��TA
N�R��p:���9�=���Đ��<��O�m J��t��z3�[j ��,�"t�.����9��}H��@XU��5vX��J�h}��0T����ُH�j@{���Fv��e�<������_��E�Ed�p����UZeF�O"�n��󑖢X�4����xf����Daܟ��5�{>��]_��P�ߙ/��L������w��&�DY�5��9,}���ea���e%B��hГ�R�(��.�����E�>mzl��q�Hǲ��c�\%�)�Y.�;��Q�@`٤�����g*l������cG�̥\Yo�J�BX�*"����\c�y�J��̩6�QP �Aу/��HL_��v�5����B߽?<h�OF�%�r�6�-�Z�Y�vS����b��c`��M��v��D�6G���&l�7�v�n�Kc!�'���b������d
�>rv���CJ�&S���F���cU�H�FkL��+ 7���DL:4o�5��@�9!}c�e�-�=��\7#K��[%xrT���As"������3�Dҕ�Qe�/�!�l]Dg�	6�a���l�.�ֳ��$
��c��D���ר��>�;�_ꏊ�azo}˻r� K�9��P�#��.�9��]��� ɨUT���E\7,��0�s���"����T���-�3�q�>�P�a,N��_���������`��ʨ���UL�9�G�%ׄuS6��}]f���ڽ��E4TP�̩�%�g;I�|�,O�ٴ>*|o6� K$�ۈq�zJp@��������Fۮ>2�i�ު�s��mD1Y�S��?�=��DCƪ�ݭ��R�(f��5����È�B�^GH��:za��c��������)��-y��|73�?�~��V;���8����w�c,�
��GE(f�}�mmƠ�F?�����VV��o�GD5�B�^�#�)�9x�]B��2�fF�7��3����2ۑ������~�T���� ��|�l�r-��ibLKAB�Qa�n��y"q=����Z���]�S�w�=����]�����
z� e#T�+�I����i�nQP��X'cQ�b��� �x*4VůQw�Z�;=�X._uV��:Ot& )�#,%-<�-��E���-��`؅o��|�v�c
��Q�"�C��L�r1O)���{�b��?�80��5�X0>>�ҹ�B`�8���+O����� Q��"�S��M�.˽�\�&7��/k��r��N:�D:�g*��������G�?��(��ب(�33N+ԁr"z�AE�8Q�/��R�����"�S��N&�"�,xG���U'�����ѝ�Q'����To��5 ��Kt�I�Ѩ`+���숲�4~Xh$"-�P�����"ßL���S��D�#���s���L/����,� �-ޞ{��a��� �r��T#��-S �]mr'�;�P"�`�v��uV4c����f�� �u��پ)��-��̤���X}a9F�����u0�|�C���$�3 ��fE�rכ(���s�߶l]�ݞ���=�,��@��.��;&�'#vR<����`j#<�3݌����.�B����e%n��u
$bA�۪h��W�o�t�!-���Q
�G�4V��J�̧P�6:h"T�M,ck�J7����[���J�N�M��]�wա`�	uI{��!�����R����˿������a�I�j���(��בX���d7���� ��O�ڭ�5���}��z���Zy�.-CÎe;�%I��oU��2FƜ��6I�q�xC.;�ұ������B���� �Z��6g���R#R���!�8���p.cD���ԇ9��G�ؚa]f�qIɓ$Mt���v��-Y�$1�,�j�W:U����n�+ �J�}Ӫ�	����9���`�З�����dw��}iW��n�E�.������*��8`nc���G�Љ�7�K5�S�L�|s��ݜv�(�h��F͏�pm6.N�B�� !������p�����Ż�k'*����D��%z�r�><5��d�O��ƭ�"�t�jنW R�Z>4�W�JG?��\'
[����Rӯ��Y�B�^�����NN��z�>� X�ܛ�@+���)�Ӭ����)B^ңnB2[��0e�: �}��-��=�	�Nf/z