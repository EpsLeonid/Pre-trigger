XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=	��%��䥃�`¨z,a�Zm��biS8����,L��Ή9���ՀMh��g�"$v��J�:�gl P�f��Q?�J������˿Bͼ�k��ʌ�5Pn�ϋ��/ZV�j�k;�E�'����X9y]�u2�p�W��}�A�WO���F{g�[~ �f��4N�.� k��侂�x�Y�El
n�5�rhD���kW��T��kA*�&�~�)r�WU]��!L�:WA���! D�)s���az�qRQ��~S֞�kK����Vf�3;dr�_0A<���ۙq$��H<ʪ !��hi/�� ���������K#ԹJ�orm����!�R;���"LL��-j�~���0�# J�4Q?!�֋��X6�� 2k�XOB�{�P��}ūy?\�w�B1���E9x�6������Y����]�|
C��.�׵� �A�2罺�P�go�%`�9�s�,-�*G�5�P���d���x�:�ܞ�x��7>M#:����8A��G-@�$y�$�����[�_fu�u��u��U�Qz}׸hܜ5�^��F�>�9$�%ע�N�>���X����r��/�Ts,��X��^m�[�M�R����[Sw%�΁�J|NC����"�\��C���~�3�ՉT�G$���BH���x/��bx!&�6=�E��O����qi���ݴ�O|�=tİ\Cѥex&�g�po�M�B�<d�R�Ϥ1h�|��Dȏ����T�����L��c��XlxVHYEB    3e0e    11505`�R�Rܥ�}D8�T�������e//fjr����eYD��Yz�M��2���X�TF�-�KkJ��N {�H%�}�k���XZaf��:����Ŝ��![� ��K���R%j!2#vs;瓎��Ÿ^J:�e�z]Mb�� �P_�[�K�Я��K���{���;%K�0?��w�VZ��W���:�Ro��'�7/�����g,���䱵��e�:����;��c���D�}%��L�RYc��8<�/n4+���R��B�F3���BL!x���	�I�9in$��:V.�/�!VAX��}Q��l��qN+�Y���ݥ
��"�Q�bjמSd�k7�"C'��u���*͵�jcړ+��q�`vOVwWs�����	�?�6B{j�)f���k�'���CO�O�h����t$���C��B�m��|Ր���w�w(a�@峝����L�?K?�&���Q��S��K�bs�o��k�|�͐	XvQ�#���xY'?r��+V:|����?��F���)2�\qE���t���mR�r�Q�bB�X��7jOn�"(�d�d.UU���*L���0��0�~y�Lh��s����Y�<�Uz���.�O�ݔspB�d��N���E��wzwa2Ż!4#��T�:�2��9L���7�+�N�s&���x�߾}����%2Sp܀Ϸ Q��C@��yBt�ё��P�pm:WG��_�Y$����t���Ƹ�H;��6�]�ۙ�<��I�N�$Grt���2�r�KB��Q��H4`,�hSg����k0l��M%׉d�
�������@��~u=(�ar�'O7���c)�.]�~<otp�BeHr���ڍ��(� h��@-�M�:��g8�oi�����U�Q��L,���@mbk��8�]����+�7!�ō�/��ǧ^�ү�P��Vv^PB\#���J�kz��̝���s�)�?O���l�nH҄7�?؎V�s�����b���<m����$g�[^ND��2�vQ���då�)�;���snj�\|�X�Vc��w��=�K�{�Mܱӣjxǆ02�6������T~i�t��%d��H��}~c�j�U�\h��y�gX�jv��J����Eѩ��C�4���e���·h��_FΜ�>���V>I 6�&�<#-��
ǩS$��(ld�A�������~XB����4`,�=t���ۨ�A{� qFb菰^:6����a�;q�㾏�꾤}j������W�s��f�ܪ��{0R��t�8�����(��l������_v�tGq��:w~�jAJpX�B�.D6C�����i�_{@	�����Wϑ�CE�$<o�+��!��k��3���@A3Y�GP�,E�Y)��{��MT�&��'-�������zK�n��g��bPb/�i��H ϛz��*����b��45�FY�?�:����(Y2�X�B�'�T��<�Ly;H�e�_d��{BQ��}� ��G��(��va�Ẋk���^,���Әz�(��|�B���z#�h�M�#j��:r���P��:Pϫ��>�A���
��.���$FQs`5ĳmmCTgi��+"t���E�yJ8�h��rv������E�
���O�R�g��>�F���!��C� &��C�R�p��L�1���Od���V�Y���=,n�~]�I_1aw/��ŋ��fH��|8�+�и���Z�^��}�߮ ��b0v��s��"}\e�<�C�+/H���@N��b����S�E��8Xе��߲d�3T�fj谹U��U�e��kW�E�P��]���6�V��jk���?0���AbRC"�l���\�2+�s��f���� kʳd�!vpNzHY��$d��vQl6u�D�kq`e� �Jdd.ĺ4xY��O���/y�`��,�q@�T��D́���R)��8J߉鈅�q�<(,EB怊ܑ+�B>9����W�o�%�ڞ)&}���z\l�d�|)�EKUp�6��@~�\�ރ����h�s�f���:��<j��=���~uF�{Ɲ�lĮ�^oS�h� ���;I
u�5�f����:8[m=�,O��Z��T?��
8�`�S���[:���ґ����0�t�����"k�l�L�����|�&DW�]�/������}4�����(�r�C�"i���TUk��;����}��{���C����s����<���u�eB��9�.^^��ڥnNzW�+u��.ll��e�Y@��z'�9��Z��ݒ�������`7�����M��M�ˮ�2,��3��5�.Yѩ�Z��c�t�/�F�t:Qd�R[͝_�a��`b��.u~=W�r#��v{P6Ⱦ�����|R�<����S���}kVo��8�-ɨ����	��狒CP���ϕt�-^"�V�Cf�Q�5>U����[���������X��t��{���!���<eP[-����!4�cq�ǲ�f�B��0�8�x㻗X#f
�uv�u���uđ�ċ!~S$�iG�^A�/��N
xy�"#lH\a�FK�R��(9�l�y%OƷfp�5Q����ldGD>D#�kL�[3���-��|����@�!���W�{`C�2
z�[xS�Z�=��X2)�:��~<g���~�م��.�ȱ�e.�}"4����nU�E��B�-���&YaDz�(�g��a�Nz�ϒ`��><)5�ȏ���8�Q�8��ЋT���s^���
/E�����2tH��'�8�-�N��E�VpV�ɗ���Ȑ���gɈa�7����7�R3��y���
��i�㗓���Ƅ1� Ԇ"%I%<[������h�h����V��T%���{�k��"!P<��U�Sp
+l����vk#�[Õ�Y�X����ڒA�Yͧ�޻���)q"/:$�3�D�%���'	�+�a����}ȡ\�����L"� �a���ƻ�?�4o�PS}�I�����3���y�h�"�����Xa�E���7��q���� �e��J�:��`jj���:Fq�Z͒,R�7�k�������62A���i�{�L7���PL�-���>�~����Õ}o=r�E mס��Vuۙ�h��~����L��׼�&�E�p�+��B��� ?P�%��i&�\��R��2>�vr��h�p�2�q����.�^�k��4��&�n��C�T�$ �֥��A��0X�.�\x����</TZ?k��/� ��|�6����h����Ƽ^fΔA��%|N�F��D-)���q��GI�9#�����Wr�8h5��z�Jhr[�1{_�Nͷ��qu�)�ߗl��+h��ta`��aJa\��?s�+���1wq�J���~B������2� �.��д��Gu��g��[㮢[�Ş�­���z���F�� ����K�܎-;�X]���M7�@h��З�Ħz0Vjv��3�A�f��Ƀ����yƠq_}[?e�!$�Z1U2"ߖ�T˂�v���|�,��2��W��i�t�Z�L��0�uyT�b�L�E5ہ�Y�� �84Ll!QM��������z��g�'8t�6c�}Ow;��C=Ր�B��4���K��M���=X#�]��\�i��93�iTP���'�)�E�H#�Nࢣaف}t�8�2
�{���[���U�(�?:	  ��g�~�e'`l�� �QA# {�Z��ώ/B4o��%h� ��Uť�^R�~�}����
C6�'��ɺ?�g�����ۓwkF�g+�R8*/F����p��"�\ ��R� �?n���X+�m�i#��j�O����pfO#1��lB��o�a�ʈ�PK3?��z-�;)���̄�8�-X�YE��#4�_�B�݉@�{4X]����3-oLF�ᐕ�_�]��k�ͼ��"m��$����%�!�$�l���������{�t�i=�	�hD���F�)KE*V�Uh�W��y7��BޭS�Gn���{���h�[�V�~��0�Q���2�h�ݭ���o7�x9��]�J�ʀ�L���'��1%����5�]ֳ��.#r�SX~@�2�5��ӭx��XsD�kʉF�5fxOT&�aѺR2[��gQj��Giss,���c���H�d�$s��2�Q}(Y�����~�L�g�����,���g��<'�3��<+�-������N��K��^�[��t�D4
�{��GRG�9���-���]q�C��:�~����J�F^�}3&�]�)jg�.i,w�0���|���w��r��ٞkN0(�c��?P.�"�z�q�d��𡊀�]rA���ÝZ]�@9n�}d�O9��\��JyQ�)�