XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����n)-���!�9��d�Q ��d���)kڧMtZ��w%L����5#q���8)&��0���cs��E%���$3ĮP �Q��;P>�qB�գ�M!�xRR]Z?Rxv�e
]L�D`���R@�"ٸ�* "�**�b.���CsI�(��S�c9���\m9��o�O{�kf������W�'B-@�s�ͼ���su��3H�_������|t�I3�)�rІ��Y�����s�5��̭�W�G��5�	�#�ˉ&Ӣ�*��J[n�h�DS��'�rH	�O3����v�T��ԟ��%��X��(ȶ���-�\��rn���^�g���.]aߴ`A���m��y�!��<R��D����� z_�ͷ�\M���Q5�<��[F��\�'��2�������}N�I�$u6��|�.9���"[*L(N���&��.��-\"Z���r�����I7r`3ň���Ct���T������`�(Be��7���v�?�4x��LW�{{����/W�&�0��-h���
����޳�y߀p�C��o�'p���E+��؛��%y��2MdbM6�D�ߟ�߿��
��a�͕��>h0��/cy'v�����(��6���6̍�4�� ��'>E2Cr�N�����fO�i#���=�D� t�%�ѩ{U����-�/Ӎ���������Q �F�-{�@������Z�hƎ^<�0����և?[��<������XlxVHYEB    5fd1    1710vI7q���2@��,��=!I�/O��Z���m���Ȱ�D=�@
�1H�^���<�?��� ��!����se9����g����iW�h�������@�cK�.����b Vm_ H\��l��<~�����3X�b߷�d�\U��c�v1��M�4�7UV��� ���e��H#d�3�
	0�jb�,�YB$�_�?!#=Db��" ��u��:3"���̂&v��2�>vBJ*(ݤ��Y�{f�P�]Eۜ[<�~�M��P��峯���,އ�Z]H3O��,:<.�ʧ|��u\���o"n	���٥A��1l- ��9��Ȇ�Z0��%n�ܣ���IH����i��c�&�X�˚�ڄ=J�H��ޒ���n��������v���c�������w��a�ȗ�Z��{"Vɱ��,^�	��,,�R3&���~�o� �F���Җdv�u��˻9����g[we,yg�S�LO0~�Թ�J���>��Xi�-M��?��Sټ�ZH�)�C��n�\aj���Tl����'Ҙ��J@�>���3�U�Ջ�`s,���m|>g�#.ff̩�;����Ճ/��ix+�d�!���~}��(�vA�\�������M!%��$@ZM8.u�O\҈��� f���<�l�a1d��ح�u0�l�]��HIRx�ﶊa3Ύ��|����B����Y=9-Ф���W�Pa�IG���t������*c�������Ҩ�������UK�fbz|���+!� !U�2�t$�g_n�F�]9E;#��t�Y�^���FTl�����ɾ��zԋ����0�J���+�7��wy�\�ʰ΋q2@�W���=g�����>PR���\}���ޗTDcϥD����B	�ɜ��~�99�VSr ���3��_�?vBG�@��^���"�wJ�X6��:��u;���s�g����Ǜ%��ܱPWy���U�{��9<��=�$�-̀u�/���s<q΃QW��AԺ�*[W&���{��ӵ�ě_4
 뎎�YMS���Or�sUZ8��y�ǅ��'�;�o�,�YJz��T]C����"��sKȓ'����T�E	3�t�Ds�W_��~�������P}s ��u`�&F;� ��<��'"���ʸ2�d ��p�Z�35Yv���/$$�Zۨ�,'x�g���W�p$�[ىX�w��Id�P?��L��՗�e�w|��e�|k�G=O!�;%
!v�n�B�Hd6����A*M:�K?ц�p�m�w�(AL��)]e�Z(�.M��Oi����f'A�C#j��-������i���1{���^�~љ1�Jx�+���iP���|{o����U'ZRzN����X�6G ��� P�D����p���|Fcq�r��~��%�p�b��7�;̖8@U@�l��j�%uf_��Z�)�(�am7�1nA�F�j#���[U�5	&΁��?��5sSS�d�??P���I�/񷉚;<��}�I��ׅA�D/�<�����`�Qb���f�WD��gޖc�n��2��L�]����p�9�?4�`/�b#��!�զn0�N]jR,�f��Y�W�5��l0���?(�>6�#B���Q��V��IoYkzH���dJ���(l���UŬ!�E�>��'�R^��Ei���rW�)��\� �"�m�}�hؿMi
}3�	�
���ڥ�Np4�0��
�p�k��3�R|� zaq�B�i�J�n���<V	�c�X��5�L.,�!��L�=��g����� �`�ɍ�0^��*��M~�:!2۝J���Cxm��>�$�����`J���-{�͇YƁ�K��1�T���4��3մ���6��_�|���k�-�c������b�%�E7��y���4���+ ���:�\0wM��G;����F�j�5M��P�k��W���w4vê�8�e���w~گB�fn�U"�}s���<��vn����?������A�[+���<ί��P�ivvki���D���y��v����xST�	���E�KQ��6��D�y@�r�"7����u�!)'�i�JV�H�dv��OI<� 9ؚ\�?�l+0 ڷ�l5z@ß�B=����v-��}J �;����U��K�;)S[�e�_؋K=Xs.u�2�Z:G�}*���(�c"9��I5��0X6B������u��'�ſ_�r��،���:��\�=�n'}��u�j �8jY�7w
��A��a�����T�����6tW��R&���|eㆇ�����k�ǔ
^���c=�;d��C��lS)�i�P8)�c>tyۻ�e*��d� o��5ĝ+n`HY��m�����5N^:e�$�v�e�8E��r9TD9K��pBR۝�~�;)��f=�8�(ΰ<���0`_��Su
�|�81ꓒxR՛�N�+ �X�ܻt�)S1f���ԮZC���j���e�M�g+/.�l���,?��5�}�M�N��T����%}$����S�Ouȅ��.4sc_*��J���Jz	�9�L���2���1�ƴ���뱙��3���Q&yJh����D����
�4�>�S*���Ὗ�2%��)dE�i{���� 2�wo��Z�G�T��p��%-&�m��=6vΥ�i �'�&e��^�K��D}�o;�`c����ێ��~�����]�G��� ,w��N���3X#� ~�![8����І��HLi9L��n�Ɛr���	G�yG����+�P�k����>ߋ�o�ΘnR}�}gS޷\��˖{O�ނ�b� ��昻��bf�!I+L��O�+.�;k�^&|�~�<�d2|�N��4��op�or�s>�0�9A�$�K�o-���������`4�~���L��\)+ӏ
� �ޅ��oR�����6�_�	ί�Ds��,��jN�`^6�Y)�I��f�q�Vwt�Ek:P����sd�3��Ia�2z>�3�;ݳ�����\C|�i;��=���-���Y�N@/�K�͖��2���^��珼U�ep��^F�J���R1�a�_�y�J���ۤ'>�XE/�����2���B6�~�d8�F����$�-���)�[�O	
̞��o��lB�x���|�\�Ug= E%���3���i^�D�h��u�sEd䒏->T~	Z�3L~����<@�~��0���#�@J��@a���OT��?u���x�si�w�`6'��s~�s�ĞϮ�(�㭀|H jZx����A�L��9[�����~T"V|��l����w4�^�������SQ=��f٨i)m�V*�2i��Ī�lw9������ �D6�|���ާ�.S�֬�5U���Ν�l�wt��ǽO����{=#R� 3~�I#�H���_5�z
���{�����Ӱ #��WP�\8�����O~�k�/��ă��W�)��)JR�[I����
�4ce�%VP���ضf��d����pv*�H\͒k~��_���� ���?\�xK�zn��6-��_�`�ʯϔ�ܢvYf��N�5U�R�fJJM��)��Y���>)�B�Z���tL͐q�0�j�$ˎ+f�+i���*�0$����n"�8�'�]���aMA��Fo=�׼�ｬv���q��6�&��)�-���� b��s6�0���tcIl�RUc���yR�^D���7^��-�J蟒���H��vف%)��{K �i�3S�oX8Avi�×L5.�H#ۊ����X7��ͣ�b;�b%�7����K����M��<��]�]��Ɗ^�V��Թ�1,�4Ǜ�{O:�t�PǀRI��/��^�$��ΒS������UZ�ҵ̏��Ou?F<VV�9�_:s+����V�83�Q�m{��s��e��)��x��e���W�l���_��d�"�6L��67S����
��;x���\ʵM�jH�lM�ࣝ:�S�uP�Tu�馃O]��� ����pxʟ-Q�ExZ=TPU2}$�GK�t�D�Kj�����"$	�zZ�S�ۥRx�\�1i,Aͺy�B��u�-14n5�L�.a��E�'_}���?h�bs��t�6$3��k.2�Xd�P<����t�L��>P���y�,<����.��C�_�f�2m���B�;l��]J�}����g����}�^���4���Y�f綵Ar� �8p���K?���Y���m���(R.�E=7�`vܺ��:�}����d��g�5_Jt�o]�U�#� ?��rA������_�O�t�C5M�'_�od�V=���N�i���wJ.q��4�J�0�⩺�~m�ͬ���ʴ�U6��G@���M����y�Ii�"�_��y��p�<���oa:�E0�>����^G�"��¿C�S��^�� >��Q�*�x������s(�#�i�%]��"���m�[�2	���Z�|uU��{E��:�I�	H���t��n>�L�����p�Ռ��x4O�)3�pb��<vi��p|��~�A�O�S��ˈ�1"�'ɎO�{9�׀�)��m�	�?�juc�Ǉޔo�9+�Ǟ_U��v�,
��� ��r�9��}A��ߢi�'���|A<��-�Bs��U����vB������a���b{��r�)G"L��	/���r8�I[��]q�+�\3i�;����ӬJs�.������~�H|�J�
$_���[(�+&�uݿ��2�r�Zt���Ҟ�E�s�R� i��8��Ԍ�o�֍,��[?Г�a��\)O}��j���U�iV��O� U��[�՞��B��>&���Y?�o�j�D:(�1�8�����C��LI���r'��&�Oy'�gv��m&^�*~v�a6�ү	��>K����*�5n�2��kݤ��\v�{��P1���n6�m3����U����H[�i�v>�Bfϰ	��^5�=H��/��g4s��/�	"GD�N�-Wd���j2�'��M���?�ʖ6����x�`���+��+,eG���o����UM^a+����g�ʃ]����;�����PJ�<N܁�b�й����с���Dᶳn_�װR���9�pr�_�=��@e8��f/��� ��6��'���n�Ip����1Pq�&n����U��c;e����q�#��:�fB��=R�]����T�X&�3��ǰ{���U�*��`�>؋�Z."�ؓ��X��~���ϼjl/����\ I����A�T�y�lv��fvcj_*�b��)���0����<d�b�Y�H]c����D_;�ka�h��5�Z��n��{��	aF�>,�-��u��l?�W�]���"�6���KٚN)bz�e	i�N5~���v�g���S��n��N�Q�%T$�z�{:Pܛ�(��!����7�L���E}��o�+�p7�Z2S_�Zr�^;�:c�y�v��װNhz*,���{��<P��~`&��a�w~&�&߿A�zf����#U�F&i�ޓ	�h���h��z0i���ı�g ǐ��Q���/�W���v�ot_���G�˸q(O�1���$�X}9�miY[��<��^f�I:�(�?��;/�۳�Ǥ�=!� ��)$���؅�Ƕ1�����9=p�bۡ����*9�C��ʜ�����ǼU��B8�L>𾍁&��<��^P�*�qt�%ꋀw'*�j�ԁ�
��Q�`W��w�3�� �6����OO��1�& �i���P�@���X5�Q�g��H�j���G;�����\p�]-i3�G�
�j�4:��t�5��H7$����%�