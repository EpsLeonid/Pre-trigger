XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x�&j$t/��)�e�&S�Χ*�U�%��%~}([��a|:�?Z�ޛ|��oA�Q����m�I2��Lg=�F�g��i�~oRq�|�ǿ"|7V�x�.���b�ش8�)��E�,�(��@�p	b�1�@�G��;��m�B�r1�^>Xn���y�JJ�w$���Y��x<����皬�#E����E<�o;���?2��W��'@[2�g `��?y 11���Dʧ�~gN5g95s�K�݄�$,��-������*������[�#�ᎎ��Ec���QϲY�g�Y�y�mn��ݗ
,�e��.[;b*J	f=YQ"[�lp�1��[��%�bD��0f�ܕ˒�|� �E��,:�����J��9�藞�ݕ��fR@�m��sd 6����%lD��pЄ�95��iT'���v�Xn&���#���U�������Ⳣ���r�P����Gw��[>���Y6+vu���yO"�%&b�OB�N+���S�뚫�a �q��$��D�d�"�� ������+,�@ ��j�=�u��g%�(5?�d�P�����[���'C�`Z�E��G8�r|UB볖�����R��8I���� *�7z�r;>q$PNddn�'hN�4U�.�n�ń��uB���N��Q�����5�r��%لs"�l��O�[P���h~A����@_[�g�{sv�)l�겤0��l�(���{�l�6�	���9F�x��ib���V���;.I��1XlxVHYEB    9653    1860������6������9˭��Q�����p�v]���th����Ő�:����iFt�Dok뤲���Ê
��� �&�w��8T�)ys�R/Ý����ٵ�Ϟ�ly8]�Z���,�Nۅ�B��'���:t���P �r_F�J��#"\&"Й�1
�`qŌ���/{�W�b% ��g�+޵��9���e�}����@
�������s�}��8��a]\�r27�R�9��������c��'������k��q�r��ė&��As�w��u�!o<�)�N�L	�"����b�EԒ�.��%�|>g\�UНH�a����!.=Q;D.s��
zq*J�ˡc�k䜱H�lCFkن�w[��J�&<�{s0Ѻ�Ty��o�;�����L��ݛ4q�˹%S��op�__z�J�,	��O}f}MW1��2�@�ґ�*s�a��$�����vHG�����gv]F������g�PDU���w��yp;�
Pu�햱5R�wn8$M���k�P;��Mi*���s��H8�?�5�R!ܤWM:�׿a6[e�,)8[�D����~��;bS��>}��W�!�������W�6U�X|�l��|�v� ����?gz�}�9�Ϛ�M�_O5�:� ����P��5u��Ouu�{�<}�d�O�l(�)�M`"D�����/�z����]�?@�Ѝ!#�%�XB�ۋ��O�DY��FNؖ �~T�@�~I&��`L�Su��P��\/vuB�V�`J�;�b�a-o
�Y9��R��lA\*��{P�5����>	���)� �l-Cj����({��(�W���e>ܺ�6*�>�33��$5�lOd;��{��l�u�Tʹ>�"k&�R�ɽ�7��3�zaD`�z��y6��ɏs)�*b8�pB�i�m�6؏���,9I*�x��Ԛ��՚�V̈��z[��`����Rj�ı/��[�KfƂ1ɎƋ�&�ݣP������y�1z�$^�t h��9�5\�c���V�gx�`6}	TvR;�ۛ�i2������kA2d'���K���TCS��Ju��J�[��p6V�w�&����%cW� �я�z\��ϠfRbxf=:D�Eu�*��`?y�r;mw ~g�bsM����9���R���o�>�����r� �wL�%����,�Q�k���P�R5oK>Q�m/>4�mG��3�ÿ��@�ʅۈql�{i���CNZοL��]n�'}���d=�g��j4	��RW��)��Xσ�-N�Q%w�CP�sw�3�Y��� �j��vX���O��n�4�̗TC���z��>T�@��4'��35�������1����&�b�2���XPL��QUVi�(�/��s"\m��;�R��3���dW�-�mˎ�kx�W��5,9wN��>o	-�a�hG̓B��(a���D�\�F
۰�S茹��|5Ҫ�E���������g�a��e�F��~	4�6s�$+�[��5H��9]"����8t���`�F�3��C�.�e����0�,�ٌ�!����U.g;��w�u�z�]F��� ������TX�5�:O����+V�����:e�u�>�����q��FJ�A�l��/!Jp;X�6��U�/mE#�Q0t�m�`�1�)�E������%���:C�<�9Mh�mC.�V��$���g�J�T�23htf�:��#�ێ��g��|�/$ r������� �yH0C�fC�=�C�KB:���w�`_���?��-I�硻�=\S)?#�������L��:Ux��������"�$�E%~s��콗U��y�@���@a<+���Z	6��.]�!���c���n
	���=��c�^�"�L��a���5���C�d+�:�"z����k,1��KE�-݈�
����9�(�t��3�Rx�@���M�:cC෷׸sȝm�"9��^�����ӊ�N�P�n�\["��jcf.%��3f"`4�i),���υ���8t~�r��?}T�p!�i����L��x� ����~"|׈1�N��{���\w��0���V#��X�հ��m��K����lJ�q�����WRE��������۴yw衣�]����j:R���C|5�9+�~zG�Ѕ�g�RJ�/ʅ�L�;=z4p|S�$ z)�� ��Z74ձ�￳
��o��?�[�T ��t8���>4n�s����3��j���V���ǐ14~�v��4�VF�z�W��](\@g��2����~��Y!����J��q��+��t�^��=�`��87�6����s[<��dI.�i����$��ڙ5��E�VJ���u�Ȃ`X��O*�H[��<�}�D��,��-\�M���t��	uun��͚Mp�h�Q�r@�7G�
�_ls�EK������P�x��R�ck:�i�#\�����%i:�=�"Y%"EjmK~�s�ٔ,FȊ��?Ď��KX��s
��4���E�SN������h*�
X?�^~ܢG�E>y�w�{$�	��:�P� ��R�Р�R^�7�" ��[��g��2 %����!;�\�(ϰ-)�.*0+���7�	�X|L��j��\8��Am̼�֥$���x��R��4j�g7�EV�r�e+F �l�1�w��uV�}�HPו�!E6�xo),y��>���r�yF��i�Ek���$'�h�1g��7b�4�����*��O�س�vi��q����gSKh���볥�Q�����;j�N�4�AcN7�^U�|�J5��I=A�XӗLR���'9@L�m��C�FБ��
���)�؂��Ť���q���jI�����wJuٍ۶��u�z}���{���2�j�Ip���^����O���rê���3B�KO�:Ë�f�U���p�[���r���f���ķF��
=������0@fo�o��D*A(�d����Ϙ�����4���y��`+E�P�K������ :�h{ʚl`^��4��E��26]���s�&�zZ���cI�#gJ3zW��/�J�v�� 쎧��*G�BךUV�%��A����� ]��g�" ^ȓ�R>�"ce�ȃ%�)�L�&��b�Ym���n?��V�
�#-IT���OK����2��3�1BU��P3���/%���;X���0~��3c5ŹQ>ӱ�S59
Oa+	W�la�˅�s�jз̅��|ȧ���M�k.f��˲�}$���WX�l֘����$Ԑ�X;7tU��TK�\��1�
�`%�⇧���޺
�d2N�C/C1Lk�y�F�zK^%hӗ�I@�W���������i_~�V��w��G�~��Y>y�x�2�	�h9�=ʴ���9����;��q�Y^�M$ $��#I�=2�r�U���kR���z7���S�y����D���.�����1G��]F�e҈S,�A��(���%���#y|)�
(�)�Bg����n��-~��X�H�(1@���T�.�Փ��K��E���v+�E�gzz�#y��,Bs��V����:��隟�xw �P�#q��3��8�?�ƣ
�^ad�2F
ǯ��v����kH}7��r9�䎠<��=�7F;Ԙ0nѬ�-�!$񝴈r�'>q@'6`�1T�ȓ��6Tإ|À[ �ˮ��z���%���ԋ*��Y��������Kqt{h
��Z�'�~-��ozh���O"��N/x0�/U�HA���P�E�2�1)��0�|z��m��a��z��y_��d��K��R��p�{��IҴ�p/wc�2,��90�����m�I�n���H�ux(l��H(:Ǻ#���|�1>��<�h"��\J�M^�͚�k,���o� K��V9�끪泫�Y��խ{�hF��2ߐ�3��G�ֽ7{�|�"����������䲲�B �9��4!-+������"��C����VaW�( �A�v|;b!�J}��ZE��Q�M�͞R<�˗L�]s�	]��v<RA���B�;�$�}�����)��Fܿ��?8&M������m�>�6P*NG�����X�~��t̩�w,FԲ�0f���5f�e��3}&'"��\��I���`���b%�
�@�ok   >�Yd�@y)b��W���ʘQ��+��q��i�뤑��bJ� �
x��F�	�X���#�w�%^�+r:6V�ab��*�����%��d����w)w�Y$�@E�T�o���1���@p��Z0v��濓�Ot�>�����ߪ��\�	���IV��N�8�*"gkJ	�)���6�􉁦��l��d��`Y�{���e
'���$��x���fh|aBceGt�V����Ѣ���	�7�BYYmnx�ؐir�������<�o�.���2��oeO�V����.�����,�h��t�}d�$��&Op	�6d��=j���!b��&��س��a$rf�>;�䵥�\���>�J�/�1+��7�>�5��%L�-6{� ��'�E�\c"!��G��B }��v���6�p~Z�+Nlj�1A�,���G(��b��b��=�=h�����}�:�ܪW1~Y�uvf��|��;��>�#����b��Q�=�;~�\.bk[UQ7��f�~a��~��'����EdfC��cJ��$� ���p`�G�Kq�7�9�F�D�9x7�Z��v�\�K��"�Y1�A3���:��1
?k ��2y�����М�>�z�j�^�s�臘�M���tZj�B����Љ�l}�p(��ȱP�"|��@mg��ʝ36XJ;؞��HwR�/��RDF�@���:M�M^�'�>�0p����Fj(o���s����l�	v� ��� CR!����k��q�NΌn�C���HW�R������:[�>�OSq��˪�3���Q�[��`-��6�����2�ߌ�-��R���\��&�:r%�_"LT.�+�B~a�����$����hd����֛^~C�ؼߌS� k�F�~�ś����+�Ah���K��a�]@�:5y�����2#e��Ԓ��Ic��a����|�:�]�o�d��H�R�%^��8�1ؠ*�q�.�$/�
�V�{��o��T��Iu2�5Ս�7q�	0��qyd�����_�ŀN	��֮�L��1���(�H���}��_�lL�>WX69�׋��0V�����e��&�(�3�d��wG��M�H�H���v�q�(�g�{���b��]��z�Y(^��8��Z;�:������'�C�R��5UG�ŌJ���3+_I�%.˸��������$81��T�e��lz}f9۟>'2��jT�́��2=�ġ�k�[ 9跭��|3=��m��*Y:{�)
ƿ�$yת.a�|�9��~���#�R55S�$^`��a�7>�QɆ������L�[�4)'��Z�5rF�ڶֱ떤ʉV� �W�~�Z�`����+� U���j\>3��a%�KN��_ߓƫN%�UC�FV����rO5���C^���kj�&Jy�jX��0�ہI:�[(�B����E�[��w��ۥ��b�TI��#dk��S�K͡�\��G9H��c��6T��A�2Xf��"��Y�,l�	d���'E ׌�<���0?�/m$c@�8E�,Z�m�k�Ʌ�)8<B>g�j���V6�󣿧��ӸD���L��}p�.D�?>'#��ݷ�R��;�$�:Q����<��o�x�W��h��������A-�f7ȸ�H�GI����2<΁�7o�'����i~i��@�Q- ���'x8۽�[}]�4寜����D=J�pը+��5����UgJ��f�8��cTb��h3�)�/`;vَ�0aT�!��O5k�̣��*���7�o�ѨJQ �=~EM��U�J?��Ҏ��\����r6j��;g�3P��|��X"ٰ=*4	�[2�4���B�ivN�����%F�z��#��a#��l�	��J=؋v�e]TY_�eW���������z��D,�Ƽ��b� �xX��<�IA��?�x���~�Q�,�j�Dk�We��Ρ���Q���䷪	��ƝU���D�@��