XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ў��j��y4-�_�)�b��q.�!6ȢI���A����w�5k�{7����}:��/���/���g��ff �o�Ά�3w�2��H8�ݲ��F1
�pp�LqqD��t���Z��j�q���F�Z<~��D�N�qMZ���b�Ђ�aG�Y���y{/����]��g��b"�38q�!co�Ap�E�*V��Q��w��6�Ԅu��Ĩ����\; ��w��f���e0� $ג�'(��!��1�Co��\���ᯆ��&'v]ypj��/�}�9� �J�14]�#"�E��<��" �d�܂V@�7M��oQ
�D��x-�п��SQ�u9Xr�&�mz(�dؗ���^A
�yK~T  )x�1�:������N�	�h`�a� f���R�*�Ѣ�W�N�$zRh�A�(ZB<� �'_�~��ñ��&Q�m��fvD s�G�)=���4-���VǞ?h��z��G�v8jm�����|�K_Y';G.�w�7X���&+:�p"����[J�&cF�
�.��k�e�0D��p�p�4#�����|1�LڇR��Xתvl�m��
�-�U���2�;��zj�w`�#$EnSAJ����֝O-
�|˝w�G���Q ߪT#��w�
�m�q@�ڥ������$����F��J��M���O��$�]���?+���E��I�r�9���_����;�n�G���3�o�L����LI5�-�Ss��.�U��PFӶXlxVHYEB    1017     680a�W����C3[�9d��J����\�V�^�\F�S�G=�I��I�rX���7r�\�n�s��<�~�\�x��5>�;m����͎�Tް��bu�����G�
���ߺ=J�0�.�\jNHƞTy|)��$c̼��tW������~�X"�i2{d�zY��?G� ���	��V�R-����!Q�	8��u0>qޖ�:��X�����ќ��S#(� ��"1`��L��G��f�6#��K5
i!D��75�?1;�o�h<��o�e)�ؾ�Fh���7���<m�7��o�Kޘ���YT}��]�F��s~�5u%aj�Z�K�b���5��S���n'��.s)`�f��1u2��7q,�ŀeܯnҊ7mb���1 <�~�����ttܪۙ��g"��Fx�X�5"��o�b�Uq
��?"+��^���H�	��$&��ш8�ş��TnUxu�f��e��~|z7*�7"��c�Ǚ_��[�p5j���Z��|���h��!��亽����T[�9��w$�?fDP�/��-YM=�����fKD�՗�t;�kX���W1�x��y�3f�{Է��=���|Ȑԏs���=���h��y���~+��})|���̼_M�-�&���0Y}ZX6�W��_b���yH͜��p00&���vY�ĵ/�E/�̱�_��4ҵ�v���,>�Ά�K?����}��F�7�=��vK���%��l<�̡$��� x�g�trN�<����p�����P���6s]e%�/��Ar�޲������]��,�M$B���5s�k�&���� (W��7FP	p���v@k�{.���"��`%������l���__����~�~�HռU^�!V*�o���9'<���ؘ�/q���	p�����s�۷;)�m`�j_�E�İ��xu�_=E�B^8���PM�1H��D8=�F����=�g�Q�������D�����s�)z�{yL��+͍����x�s���7H,��\��7��`���l�E/̒�ӜZ�fS�-ž�N���6��%PV��b���^����6��wa�A��T��'�k��J��TD��-��嚎99��5��k����aT��V�	��}�Ak��(�$�?I�p)��(��M����M^eF�XwR&wŕ"\�f1�м�2SU-�V��8��Zf?��^0���X�gv�F%vG�^�9w��*K�S ���K}c-�
@Y���0L&Bӿ[>�:��G��yID�o#V%uJr�Ln0�����0nZ����B�Q�����M���`*�jKb���W��6�vzQa+Z-).��J�������y���wol�T��kд4
Kc�, r����]T�Xi_�WbeNz�����*��}���K]}����:���v�9�s�qۙc0f��V!�s��}�Qo��d��;AW���ᾊU�)Y�P���u�����琻���2���������q�Z���yk-F�w�M���!����&�T�C����cI��&�,-вO�e�����
+��5}��5L�U��k�hg���H�AwLf��1|,�`A����1��!��gA[v$�!#+