XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����&u���O���t�	�����������w
��m���̜"5�0�L�CJ�ϕ������W[A���O����-я��б�w�Wӻ��|�~I~eǽfů7 1�C�q�ǌ��ܘ�m��н���U��,��8�ө{�Y&i�9R�.����-;��(Ŗ��s)F�Uf�n]Z�jc0��C_�{�B/^���蝖h�"M ͭ=���;�j�z`9V�A���uB�5���sӋ(�Kc�|~�0>H�	s��MZ>Q���Ү�L�J�hɏ��B@L��j�!#��ҩ{ c!|���i���xq�t�$Y��Y�1{g���6�:�"�����k�;Ca?y�-$�( q��u;	r�V^�UӰ��>��[�-h�"A��[OA�!h6Zz7��X���e��v�J�,\�;��]~[[��(��J�μ�{Rc�.�85�cW�
�\�W�P+���2��,tM�V��ۜ��|�-�'gϾ�2z2��1�0k��%೷*0��+�f��x�0��iB�TXg���eS�9�)���P|,Ct����o��Dm��*��zW��b�+gC���}�Ѵ�v�+P��	��J-n|�S���w
�K2Y� 'H/�;Ң�7eY����ǅ�T	��&��^��q���~���i�);1��%�"�
7E7��aFN+��TxF������P�m1��\�����pjfo��wB���Ĥ��[\
?.�{�o���df�ɀ��8?�瞡���!�_ u�� A�XlxVHYEB    1661     760���T���r�M︦Tc�E�;`�5�+)�D�~�ht �Y&U�<�la���X��iAwȧo	�@'L%GL��'�>���s��T̡�pe�ѧ�S�����i�|5�6�ܢ|x��-��L��R��RRm8�IZN-)-�K1��Xn�]a�� 7��j������%U7�"����m ֏zO���Ɋ�a�$44�H��":��ka,g��L�~�a*���Q�.ϳ�p�1a��n�:����-g�j�8��OQ�w��۴�+�Bl01=����d,^Ԋ�l��ͤ���\)o4�����&�����2�KӤ�,��m�a��`c"�U��b�0귚�T����V'I�wZ�kNkU@�(y�e�k�A� T���%�dfL|sݕ*�}�e�T�W?����݌ER@�{��_�%�%c��%I$��n%�w�0�a�#x6λ%:n�����w纊(�����1꣠a���IiT�}����Ҹ��!xS����۹Qa����(��D��rܻP`}�A�>�y�I����i*�;�F!VjČ͖C{@��:w�(���ߕql�,Vi�Bor���$��j�FU�H�"k⒱�����`9���l4HwT����P��עY��aYDj��l���B��"F��� w�hˇ+�]�'#�L�M��K�}��̑�J#���y3�2�$�lѦ�M�~�*�?|�K!=*���`YHR��B�'�@�,�\~�έ1����cW��Cە_�MX0w,�e�x{RFj��F�(Hp�_(J���7��N�S1�PL���&�['+7��[�D��ا)���i3
��=�td���R@��bM��v�76`�Q�~��hBW�i|)X�d�ɼ. ޺��>��A��SB��2vM0�5qHf�R�����-U@�s+= ����:սl� ��IK��'h��Ў�
�v�A�܉�3|���>�I4Rl`-���ȋ����j�-�'���^�+w�-����7:�����^'�Z��:&^�o̍�4W��2 ����O��1/���(���Á�.���x�Y8��4���������F-��T�����	T��"�g������ ��>�l���m/�jiZ1W����U�?�y�k�"?��������FB�}���)wo�����x��t�����ۤ��O1�W�/.�ur�0�����3�g"L�"q���=�ՁD�(���_�t��8]
�`
�[�옄������\��!�xY(�gJS�­���I5nn{�#t���c���j7�c�Ȉ�] H5�M��-���7�>3��|_q��0w��z���r���HZ��}i�Mg���Sd��K7Of�ߛV�a\.Q��d�dsܿaO4����Y���&��(㔔Q�o8��v@}��'S[�W�=[�tgW��67lB�����KY���O/T֔������6t���:@�ݺg���=<�K��F�K(�5k&J��F�Z�,Y�o�
��cd�ԷKT��uVs�����btWr��h0o��E�	�*O�N
���v�޲�hAFD�-P�ժ�iB9��U��|+n?nsNr�B;�S0E)0s�M�����L�1�HY�Out3���Kέ����ؤh<O�)a��(��,� ޯ�����|9���ޞ�����HzՕ�-�b6�8���Wl�iH7S@'s�^��Ԓ(��-B�1W�C�RB7��5@�����s�PZ������q�\<�ov~ь#H��.�Ux��+�`{L��`o���GCc�*v���<�f3� ����?X���Ң� ����+�NI�� ΡڄwY[7��oXQ4別U������_��{��������
�