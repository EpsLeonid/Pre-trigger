XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*tL^B�pL]9�1��6�F�E�������V�y��V^[��^�~�3��WUG���P^ꔇ��c��ع���3'���̆M+R�X��?�4�>wQ�T�0�FIHSa%�����֏��3_�%M��آ�>:��AQM�(w��p)�cW��Gf��|��������w�3�4�E�ikZ$$Iw��~9�O�ʫH�����ɞ?��=��"dDZ�yZ�i�����AWD%�t��J��*f���y"W����Q��u�0*g[pqpw�Ķ��1FH�sV��~�����6	�vp����ң�ͫ�\��n�N���,�A�Y)p�ᑑ	�.����_�s�^�M\����>q�)N'�R���\9�w�eQ$�`n���{��SAc�)�Y�GV����gZ����pO��ܧ������9apec��^�9m[:�&]%�˹�+��\ߏW��!3Ehv2@ⷵ�7;�'�mp�[�a��-j�1��.�{ǝ������|imu�ɷ��~�E�"��Z�0���<�ǈ�7����~�s����/<2�S���a���A���/��>�t)z�RgLu�:-��k}�Nm)ǣ�D�ߓ�`�]���Ff�HJQ ���(���q|Y�����^����p_G���J�sT`�%�X���8j�M�X���V����
�5�9�T��v��`}��� ��7L��ouQ�҅�Es����)*-�{CF#�-n� �H��3��=��q���DsF	�-�gXlxVHYEB    3292     b80>�'4� _� ��6�<�L������i��w��g�H5Ɍ_{�[��أ�X��q,N�j��Ҏ��j��3�4�����6�CsJK_@F�;�D}>�'�����1�
A�����J/�8�}��i�P�U>����<��C��_C+����K�E�"�V�4��L�0P�
Z��4�Ɛ��6���g���2HZ�읊5|��*����>��l�,n8d-f���_�!(�*2�-�`��F��07�ɲ��S��߹�f�dA155n5���#M�R�1C`*H2��c8�����5��]U��o�݄?r�;�T
��{��P�(�HE���UԮ:_3pɨU��>�w(_Q�Fm 5��>�����c�L�o�o�3����Px��؇y��aNs�]�'3�[<���Yn0#i*�h�:���2'���&���1[�jh?�cCQ�E~�^��tdԕ��:�v���}�����o�
$u-b-4	$��W�#�������\:��/��W�Eŭ����E���D9����k
��^IT�Z
�r"z���>��/Z��>��~(��V������j5�*:ȳx(��h����'o��|S@��s %l��V.@H	f
X	��8f�ˉ:G�@;�c��4���s��oha?R���>�>Kɕ_���Nm���Ң����F`�^LJ�~�?�fS��4iO����V]���ʼ�Ɂ#Ƿ���sHڲ����|}U�q`KX�ԇ�Ky�>��!X�9PS�g�.+������+z[�kJ������\�	Y����G�r=|.�t��%B�_���1:�����J|�&���^�U�@����`3���b'�E��S�w<އƮD�������W�
�Q��K�V�S ��G�P~$���3E�u醮*diS���^�k���0��B�k�w�(;B1�q ��M����,���=�?t��mql1M6�b����酔I��=;d`��vB�ѵ{|�}�'��/�<-wJ���9�GQ�ѷ�Pc�1��1������wJO7h%`а�N�,�kn$;�$�A�M��o����.��)d��k�r̅�1���e)h$]M%���9��G�̡KU-��'�(���[��Qv�e2��=y�9�X�1l+:�4��M��l�oeq�8��o����>�n��3Ϡ�)[6��j�c?���A"	�e0�����W�ߎ{,�}wcP�]}-.�sG�T�|�֑�ߏ7�8Y��"c���Xg�<�O�����ܵ�;�ږ���8?Kh#�=3f�Ip��"�f����#�v7�f�+=ȧ|&��U��|C���jڵ�5(Y}��y�/|*�R]x}2V&r�f�3+9��ЩLm��iBʵKz�w	|>Ba	�E�����必~���������~+�/���������~�����&�P��*�!���znK�:���?�s4����ň��C�+�L��	��Y�Y/Х=K^.��d����D�>l֚����5�c��Fuۏ$�3��Q=�ԂB�_����,�I��H��N|uc�>� �_qo?�ږ\��ų�C1���2�ZYq�����`]��|��?���I)��-�˭uI�4 w�(�䀶��80��-]�Q�@��L��}u�vf,�ڴC�>���2Y�E�˳������s�-��{��)L~"���gzf-2ǵ�Hh/��O�Uz��=ރq�=��5N5�Z'U�c'ZT����'0�\��+cW�kw|JL��	��|���oD��@�����v�O6k:�0�q���q����㶾����;X�����Z�h�*߆ -N%&L��0s}��/_�8�A��(���������li�#��j�Ie(!*�˄wpbuSe�Qv�N�nKt]���u��1".�-�#�J��I}���Ic���� I"�/9g��~��7���Z&YR��iP�����r�*��9��h#�fq�l����S��٬�L�Fk�!�����W���#����mrY)�KC��gTH 2�z��^n5U��6%)ɚ5�:�+
%Ca����t��)�O}�͹�sRa(��x.ϔ����Ū���y�:]�@[�AH�W�z��C6!d�}��]�W�:����0Mt�ٓ�GϪ�3�ag"�Z��^H]ŷم� ��~c�q�G7QM�U2%W��n��A)3B�z汙3�/i�
�_7'1��U �J�(�O�N��?p���mmɍ��h��I�"��}>\4:���ZnMd)HX[��Z��f3�V��6�G�|
�Dcٷ�}��&&1�S#ޜH�3N�?�CXG�*���͜� nPl�j��!�)��s6�0O�� �β5k��{ֈ��n�kd����ވnưn��1ˑIwM�+����`�l�i,���P�h_&�6/xt�#���(�]�w�x�M.{<J�E�/H��_a;���v`C�T��⑍x ��8��a��,,��y܁h�͘(`��z�l���#�ׯd� �����z�|Qrv��̈́�E�W��������6%	��� ������ܠ,�ۄ��t��z{u��4�"�V�p'�eP�="d�)GV|��=t�x��x�+RT0t <U�@ �f߭��"'ݝ���ޚs��!E�A��XOD��ih1�s��mWW�3r+�X��:�P��s����K�Y4���M�dR����
I�ޛLMC�����1	N/r-�OC
�{�e]�"NJ�Y3��IZrl-���L.8?=�H �q����,�y����h2��λO�T��Z���kH����V�����]|���W��Rn1���ܾܒ{v�c�%��f��v����dOj�b�mB�?LtZd��<~�֭��D�W�~{��q�\N�:ۭ�j֧�Ӧ