LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY system IS
PORT (
	ETH_RST_B : OUT STD_LOGIC;
	ETH_TXD : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	ETH_TX_EN : OUT STD_LOGIC;
	ETH_TX_ER : OUT STD_LOGIC;
	ETH_TX_CLK : OUT STD_LOGIC;
	ETH_RXD : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	ETH_RX_DV : IN STD_LOGIC;
	ETH_RX_ER : IN STD_LOGIC;
	ETH_RX_CLK : IN STD_LOGIC;
	ETH_MDC : OUT STD_LOGIC;
	ETH_MDIO : INOUT STD_LOGIC;
	ETH_MDINT : IN STD_LOGIC;
	CPU_JMP : IN STD_LOGIC_VECTOR(0 TO 1);
	DDR3_A : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	DDR3_BA : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
	DDR3_RAS_B : OUT STD_LOGIC;
	DDR3_CAS_B : OUT STD_LOGIC;
	DDR3_WE_B : OUT STD_LOGIC;
	DDR3_CKE : OUT STD_LOGIC;
	DDR3_CLK : OUT STD_LOGIC;
	DDR3_CLK_B : OUT STD_LOGIC;
	DDR3_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	DDR3_LDQS_P : INOUT STD_LOGIC;
	DDR3_LDQS_N : INOUT STD_LOGIC;
	DDR3_UDQS_P : INOUT STD_LOGIC;
	DDR3_UDQS_N : INOUT STD_LOGIC;
	DDR3_UDM : OUT STD_LOGIC;
	DDR3_LDM : OUT STD_LOGIC;
	DDR3_ODT : OUT STD_LOGIC;
	DDR3_RST_B : OUT STD_LOGIC;
	DDR3_RZQ : INOUT STD_LOGIC;
	DDR3_ZIO : INOUT STD_LOGIC;
	II_SPI_SCK : OUT STD_LOGIC;
	II_SPI_MISO : IN STD_LOGIC;
	II_SPI_MOSI : OUT STD_LOGIC;
	II_SPI_CS_B : OUT STD_LOGIC;
	OSC_50MHZ : IN STD_LOGIC;
	SYS_RST : IN STD_LOGIC;
	ETH_MII_TX_CLK : IN STD_LOGIC;
	CPU_LED : OUT STD_LOGIC_VECTOR(0 TO 31);
	IIC_SDA : INOUT STD_LOGIC;
	IIC_SCL : INOUT STD_LOGIC;
	mem_addr : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	mem_wdata : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	mem_rdata : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	mem_we : OUT STD_LOGIC;
	reg_we : OUT STD_LOGIC;
	reg_num : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	reg_wdata : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	reg_rdata : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	clock : IN STD_LOGIC
	);
END system;

ARCHITECTURE STRUCTURE OF system IS

BEGIN
END ARCHITECTURE STRUCTURE;
