XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���q0�G���&>d��L�_��~J�ZV��&&3(eN�Q�	6"#]4��>.���f�o��%��u�s�]���V��qh1j2���hN`��h����]��� P�M&�ؿ,m�o-�Nr8��:~.C��p��(�����gZ��(��߷�n���ځ\__L=M�Sg��Y�� ,���?�2���k�;�x�t�U�5-.��� �������T:��i���C�a�6��~�紋�#}*��颤� V����X�p�;Ǚ��I%�ɐn�ı����8U~��_��x��M\�Wsa�����@�c� �;.�͞����/�u��?�-�z�����,5%OȨ�&N��_��u0�_�Q�34(%���l9+�o(�4TšJ��4�rˑ�~�������ݣ3��gsn5������W���>5�|�ބ��tz��r�QX� �T'��d,d��fu��n��ӏd�H�A�-��U�]�r�Gxj�cZ_F9���_8�s�A��NM�d{�(��fW��KKST)��@յ)8�=(�U�+���祀��سm�d�|��_L�/y��-��彋3�;�%	"�{��|��DQN�ѧ�QgC>yRB�>�U�D��;�����uhf��|��f	�F��*Ûo�?�kb�i��qW����#�NP�OPD��*(+����!Br�˓��E�u����Bۖ�0l?ÀK�^rHڌ��ū孬N�����RR�ߑ�",�X�b���ڃ�q���j���XlxVHYEB    d81f    26f0E���uh�&��	U,�$���t9o��\k��Q�H��n�g���$�bK����?v}��F+�j�ɀ�}���.lW�vr�{+E��.YŌ�Ŷ]7����	���6j�V\�!��5�$���aQB�7�'Q���A!�7�L#�q�D�J���Yuԑ,��6��A ��㤗�g�я9����`��dμ^Jc|����G;�.mx��+�ר��y}B���������,:�Qk��	@��b�,x���6Y�{a#O]q�9�i�#��[�9���ق���1���>���gڱ['m��a�:��8�U���+��v�������Z��_��}?��5�|'�������t6�p_ �6.=w���M��l|w������-�њ)[�y�����n3�B�(S�KWb�y=�����&k��hڪ��jV���\$0J�kF��.�N��]���c�ܚ���H����H��򁠵�m�T�.5�a�#A��_;�uy!�EL���c���(�L��a8u�e \g�&LLss�w<,��x��!�v��!�=Դ�}pֆH5*�������j2�ˑ\R"��6�"��|�Y	ע�Qخ(��:�����G���'Sgl����[pJYSL�ĥ�1.����)T��{��y}��w�~[-�Ը�C��(M+ppk��w
���}l�kߝ}��<x�3��V%��#�6t�T���/����I�bxdB*8���%�@>�&H�6��0�=A\�L�q<��$Ѧ�vd��|p<��f�3���/Ȧ��eFXcFA!� �>�'���G�S�h�v��Pt,0=���t.�cx�:��&XK@��m�b"�<`}n�WP�_��]���ӕQ2W��w���{�]!o���u��kXR�Ei�e;�����c|`慮i"T��q��ć��hԨ]�d�������+��SX�ʕ���1����������RD�.V-G��2�P��ź����6d+�b��"�u^L	_�]��ē�F�Nl������51kwN�z��W�<����v�^K�(~���v��ㄼ�|�d~�w�f���-WC��o']Z��A[fL��*����DsW��\D�%�g�/~B�s��wC��rq+���ȧ�a�:!M�x�}��;�!?)�lk���oJ4*�d�375�����>�o��4k0�"�Jj�,}RiC���U��S��\����d!ڟ���,�Rz�� Bp00�ǈt	���n���i��-�!)�΁���{|o��ezɂ!����#~�肩d����=C����8�hK���u�L��ޖ�+�l�]�A7_��E���a�Uc	
�3��?���h$�O�^�ŗ���D�@4����J/;���3��}�i|PI2N�@
�a�B�OU���Nl��e�V��;|u\��#��8���:�y�H+��M���E4~�(��L�1�����L����9^fB
�E��J��>����Ҡ�Qb��j��4E_h����$����{2J�4ҋl;�� )��~ޒ_�-���`�?oxǥ�-3������h\��uw�b^8�r�Yte�q250�EE��z��NٿÐ��I��j^}K���W#TK^���	)WP�}H�PjT%�ƞ�1�.�./�Ə�b��V���n���!l���8��>�d����o�������Um��$8X�J'��c�Yx���qi�3�(���7��2I��;qQO�IVW�1��G>^n��h�x��/�;�=��(���jm�	d���6�Plr�\��`N�0���>gHZ)�-k%����Ʀ,��~B�5�20��|[[����_�;8�[�w����r�����(�����l�3�����+���J��f�E������S6z��#{?��!���\ů�G[����2"�7@U{!� Odl��ӥ�-$���(�n�m<�p5ݸ�^�<��.��DڗI��;1�z���7Ԟ���{ْ��D8�:v&�Z��E�
�K���-`F�K�� ����D�P7�6<� ���볬��'[�[%f%�1haY���o3=/��fn>U���*ai����F8V�)�u�v�H�iT8#j�z�����	���5bog)�_���%!ƣl�Xe/lx2d�	��'&�Xd0��UgىۊkcLSjh�>����l�	4���rH���mon�֍��}��#���w^��l�rέT�4��I����"�R�W��!���� �b�Wt( ^�0x��K�I�\6Q�Ctr��WN5�P ��ۃ���q��?!Nw�?��%��يc�R��{<J�́�ʹ��@�٬ȏ�q0��1�!2{\r�������*�~H"	T }U3/y�+މcwcn�v�6�������+��ؓ�j�	�����%�T����M. /M��hO��N��wgp(�+�\˖��uz��N�؅��'�49P�`+�	%տ�~w�l����TA���!=XD�P+��'�R�g׬pAw�E����<��pr* �9�?D���A�e1��sj���s�|�I���ׂ�[�UGH�׏�:ع��P�w�5o�!���)�g�4�a���4+A~����.����?6�F�"̻�V�s.�<fv��������,L@.�N�9���,��C]1S�+��{J�^*;�I�%� *�����~s��uZ��Wa�ޅ��Ѹ�vN�=V1ח~]=jI]�y֊��A����J����8�"h62���O%0�wKNK��lA7��G�ɿĤm�.��m��? �4����Z�o�o툁Jſ��ⵕ��#�����݇�vA���7L���&'<���O���:d���X��p\���c���j�h�:8k��s:\����=�4hj;Q,�}�G�5o���V�8��2y� ��Og�/E�
�H__�I�Q`�_tz�.�
*�R/cC{/��� ^��c�E�Ʈ�t �K����������f�����=)�^-U�����<p��R�����M���߀����G�k�,����-�T=�u���c�?���'qz2��}���᱄��$��e�ZB|�,�����z���>���qt;�tu+@H�'�➊d�G���"�NR��ܳ%�`(����B�Ԟ	����t��M�������B��1R�L�<�5�x=�M�H�g/S"���F��>�MӨ�-��!�\:����^o�,=H`?�ʛ=s�~�;2���L���Y�����
p�6q�a���\���0+�.����J_�os[�֮��B���3�`ש	xK�H�-w���� �ΤO��C�1�r��[�2j�>�=(������)��g)���Zm�:Y������8��HW3n
���R����cr<��@��tPO�'݋�E@�t6F�rU.�I^���I^N�N��#� �E/�S��!I�+��Q������^Ҿ��Q�����"�J�H�$(�3dΐ5H#��|&�Ӻ�.MX�P7 �s�q�*���̴���OV��M$���j_�@|�Zf_Q>^�/W��t��^��$�d��A�d�FP����'��B��8��([P���䞆;g�	�7+�h��a��ny0&]�Wg�����JD  Z�mz��ryC�.W��w3y/5Op�=��	�Ö�22�j���N�����]�O2�XKҋ�����;���D`\��_Ic4�A��FQf�P"��F�gY y4��z�4���I�i6��zs�����b�;z�&'x���ɪ�!F�п�?Y�W2L��G��t4�A�^q�
�n�Ns_�Dqn����h�BIiE1Hr��T�k�\
w���I��0��Z�� ��voSVM7�Dц�cR�Ɉʺ���߬W@�v.wz'�=�HO�Mi5�/Ĝ��E�D����ả�����W�bIS�׌����:�&Mo��"t�І�ُ��s���e�
jnY�$m��%�5�x�������&�~��K����w�#��7_%�ʭ�<�v(l5�`u(�C{8F��r�^��H
I����J���P�,aߍGq�L�F �u��=�e�g�9�~��*��qT�7G�ė���f�u��k_���٠K2C@��Y�CP�jRNg��k�I��YW9}V�*����=9����Fw�\R�#s�?��̺R�k��6���Ȃ>�֮���=�P2�A�y����c�w��j��oj��UU��ʞ��'�3z,�.��||pC�/mEB f��,݊J���$f�4�꘷r�fȗ���h>���ȵ�����CZ��dn����L��\���b��:=�l����o��_߀��IM�Q�ZQ~��3�L
�"�2$+J�q�p�1����ZT�b-5�h���FO�Lj)�Z�b=D2��|y7��0����0�I�.ۘ��	Ns�vB7&�\X����5��*R�C��^{����޶屘71�͆D��=0����ejh3���k�7�\K�#3�\��`��G��� ?��U�X��y֢ ��Gk���%ɶ�h
?	=�9�e�К����JF�Ӛύ��;4Ǐ?u�Y�2>��������~�i�0(!	8�u�6��^�@�7�탢|Rg�� �+��;���N� ������!Me=*[̊�c+fh��EC�S��2�W&�@@�5���ZúPU��E�'|5,���˪ؽ)���2H�s�f1�IRnn(/��z�a�[mU+��������:N��(/�����ЎU����R$�@H1�5��Uun`XI��WYN]�'�ނ,�f�` �R3�
������]\,����;�T����.��8�1+�g1>0�*qc]�,���S���eS*�-�Cl��
��-�v��V��_����:�^�~���3�;�47�ed��M��[M��E���	��H�����:� v��}�@0�Mٗ'|�דA���V988V��"���'�
Ӽ�dFW��؝�Đ}pɭ,�/߾��'��=H��9�mA��G)��I��E?���)��׻�"#J�x�+n�#m��q�j�)��i�X��a����Hߍ��MKx""m�@�c���Y�-��97�)W 2Z�Y0��a�{^�4���f�;�x�bJ��+'��@�x���㽾��mk��	gI�_�Xf;�!K����Kl�(&���Dt�A�A{֐�����~}<�B����.:J"&�ӱ���?��P(����@��N���u��ź���9�'IH�ƽ}�S��ovrt����f������T�FgU(�IX�A���_�I�I����[ʘ9�z�7��0��qK�j��a^��%Q��%�LH���X�sߤ!����7��k���Ϧn�YZؔ��Q���T����K=}�u9a�GIx�C�{㓹�50}�����SD=��~�}��K��n�ʀ"�G�4��B ;�x!���&`�~��t9>��#�$�&B"1��lI�f�P{������X��M�8���?UQP�-�ʊ��럇���!�U+��>�&�}{�H2'�����}s�T.�M��n-1�x��!��:y���v�$�(AϢ�H�T��2��9�7�n�<q&�W0��W�7�,�f�rS�ۉ ř����p-]���0�qy��[(�_�0o;�%3��;�^���y�9�Y��9�F���I���=i�6��R�-�ԛ���p?�Q��tM�0������?�iRߐs�
�lY�Q���@��2�LZ+ø+�������R��4�7�Ν�<Z �	�"�KDa�$��4��1�@�c�/�gXFp�87��(��;Q��@��ʐx�e����[Ud�7�&+��6׿�;b��fO��a4b�o�7�	8�)�;��
�ή�g�-�ǜ<�yΛ�*����Ci��cɏiH�{���{�O�;(F�ê�}l�R?�y����!U�mn7��kߞ�d!������E��b�c�4��P�o�#9��'��%h���^.q\�|��;��X�\]���CxSJ �M�U#?��%F:^6���-�L�[�=��i���ӭ*.�/s���g|0̧=J�2M;4��TR��S�7�M.�a��@��Z~9��V�+��ڶ5��@P��!�*@]k(��|���*miHgk6��Bi�s^5x��3�o��ڄY�/��_�!Q�'�ȸoCq-��S*��skC���HTj�J�zN��2g�t4���#�1��(�����hS����BU�]��`�n[jX(�ϱ�T��L��H�FE9��ׁ| �b�p�S��η��6��Y�O�ۤ1$փ�7d�3�M-.	XX蹑m������D�:��d9=_6�,����F�g��>A W*��D���!cJ���dt��`����$�G<��17}����P�oȲ�����)�Fŭ٦+�S	�D��"���9
�����z ����	�n\�(��$�u~ov8~e��k�y���^����R���XtT�~�5��Ps)�����"Ҩ�Й���U��`�g �g��,�Cg}�!_7S�z �2�N�,�ޥ�"�5�j��U��cWTь��/|����
���\��UW��8�b��=��?�ǠnXؤ�+DF����+]��Kt�M��B�Ð�D��v3qEFxA=�d6�!��`� ��[.g�x��j$X>�p�He�ńA����>�'��&�M��o�YC����މ�2k�)�����2��с�TU�����.��6rw��B����'B�Z)U��
7�v�8J�T}�|�����p�j�p��^�,�/N�,es�4�O��5��*�n�9����a?�ſ��?
\̭c��`�6)A�E��l���~�/���Qd
?��6���7Tͫ)៬��~vF��WC�69��-l?��R:":���
SA��Z��U��q$<K��Ju�t�4�/(�B&�h�!�����E��$	�)Ղ2O7Cry�hMW'�H�ҍ}�+� lv��P`�e앤�~!�j^�F+�KuǕUK�km���/���8����yڸ#9�o��{>�lʼ���awm��O5�`ND��?��fr�FUdqq�:�lN��$��\-!9��hzG�S�T��w�!M P̕�|L�im�AF���ב�#T(�S�4��\���)����qbS�i��'Du�z���yqT�ϓ�R�Ќ�3C��!��@:�i��]���a���zI���1F��pS�{���>������\�_o�����rxy�� :���t���nX�\V^7��yf>�]lk#���_��/�shxvl#�FZ��:�<}�!屠����1<KZM	 ��dς�ةd1��ǹC��e�#S�{|)��h))M�$4��~�_i/�'0���u����fI �֤m����<AJD�����z��Eļ�~�B�%�� ���_M1c���9�m5��i�S�K��Bg�� ��ˡ����u�t�V���o��Bp"v��s�n�,�|�s�v�e�+HN�.~!q��.��*t���l<~j�a��(Q��yi�
�<�M,�9�^A���@E��h�ο!�p�c�Wmڴm�'riz@���!��=N��=��5X�|�&���<J^/�)]YFm��B�l��&�X��@�H&��]	��h'�����>)n��r��� )�9�,0��j�P��!�l+m�Sc���~�f̑���o��ⶖ?����]���D���_Um�C�O�&ʌ��{��i�G��rmɁg臷 3��@��y�v�����P�1�v����S��L�K�NYLPs}�,mpV����f�%�O��me1�~d�,C��̐��g��;��˾����(BD��@�(K��)�.�YD5�d?��� ���Hň��p������lu̲��ʟ��Qan��8���>��g��BT삪�z���F��E��Ӹ���f��_����;��-e��Cُ/%� %������MvQs �R�X��ƾz1�X�1���ۇ��+t��ǋ�e �t�I_	�a��X�ܫ�>0`�=AK�sE�V�����h����N{ ���<㥿+�<{�*̟N��}u�u�({R�τ��qċ!`�5
!���=^��B�C&�v�Yޖ�*��e��Q�i��E�͔y��<L]�CqA�W�u�N��<b�E�>��r5�K"�����i��-ܯ�{��gD4�vH�k�?!巢�uq��@6֖7�|��k�����p5��S����5�?V]��u#d��*l���Լ��f`�����'VE�G&��S
��E���G䀘��.30�f�j �����K��,���n8��V�֧���|H���r�l���T����?����X$�����B���B�HH]��>kRg�߲-��Y1Qq��Oe�
��C��Q��5s��+��� �]7q�~�M�:m�r}V�a���=��Y �,�S{g�f�S2�o�O�.64kh$xߗxp��|���c��U_�y�6W�՟EWmzH�8�SǪm�u:m`��d4Z���E�oO�H���x��4I�ؙ�m���;����D��׆o`�rX�*���(�i��ͳ�bd���d�&$.8@�<�NR�"��-�h�� 2W]�t;�-�}�q������<�I�]D����~ڝ@�
�Yӂu��%`�����U�P�!�T�5����o�1��:[ԓWIS����!K��֚Mf�J���m�6狇INp��2�9b$�z��xJE�cUB��ί|K+��l��ׯ�BRv�1ih��E*;�{�5gSwԲ;��Jb��X4F��$)���[�^u�N�SN&�z��S1q'I*�a�́w塥L[���$
Դ��Z��\2����~(�� )��z�[�?}+�:�l�0ڌ���� XR�B�xI�C^8^�P�����f��7�[�Y�c�|�uسD�E�BbkwE�գ�p��!ŏ � G��L.uL~Eo���%�\Î��P��N�c��fJt0�V��2�χT�6��Z�vTM�}o�#&/���׳g؆r�Ou#�z_T���TAJ�����i�*S����>^>�չ���ht�|Ҳ�}��R⇜��ߖ�s.���?���s$r��}淏�.%��Z�xǞ��m��jcC�#����է�/QKMij������f���3H��z������g;z�N�k�my�dķ��,3���F���i�l]x-g��s�A�.tي�.�_����U�3���o��>M�ԩh�6�o���خ�Hp�@И���qbe��(�"��9�@��ϩ�g|�=!�[tirt���e�,�:��1V��p��yx��1�0R�f�ϒ^o�v�vm�MY��,Нu# }��u���s�V?��	�O}�����{����Mw;w\u2��Wr�-��u�R��'�T|J'�i]��"���Aw��!墺����']�j�B�L���V��^q�N�^j��J��S���� ��Z��/��<gs�l�D='�pG�Pibط #3�y� ��$���x� =��L��ߊ��]J�ܦ�р1��B��t�t�@IkɆ��`��[r�~�whv��bg�듴��}?�ÈI�@�B�7�jB�ljL-�T�o;oXR�qq}�\b2�xv*/��Z�;VK��`>���,������x]Dq�!+��B�tH�7HXSg)�|�Sj9j���p'�᭸��8�}�A���dRm��^�1�*y�t�|��a��n��A5�����sƧ�2���1��畆����?�ȣ�Ty�}ib��	I������V	�w�x�����l���f��%��s��Y-�t�"Y��wH
b~�C��