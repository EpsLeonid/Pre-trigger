XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:�Μ��l�k����oo�qq�!��)^�٤�.��,;�y�u:H�e����e(ۂ>ɾH���!�f]"ǽ��)#[$F��l�<Ѫ�I6ө�n��-J)�PW_3�M&��G�����cD�~��J���Ȕ��t9�N,R�8ŏ��-��Mje?�(�.�3�rH�d�R�7AA�i��%�Jh1�������%���!0�ąҫ*Uk��M�yG�����_f�(ة���]G��8�x����iD��̽]J�&?O=�`�Qq7O��_�9t��\�2Z��&���L��K�nH}_36?����|]^�Hv�y�9�mn��{�C�W{�,�1$�j��c�[��E)@�j!jw]��5�8��~(x�%z�K<�r)���eE���Ām�s��Z�v��F����'"�n⒴kkq#3޻������O����� �=��+����yreP(�9���j`�>SD��Ch)(�mǱ�&��n%D��Q!z��ax�@�y�5�e	PN�M�ӷ.�}��c~x#��|�40�Ƞ
6� o-�5�r�^]�pEP���M������Sgu�$I�]�H�)�Y���_�'��TY��0o��8�d{^��Q��n䅀A�p��{�b�s�;\�>Nz�{��wE�W�0h����n3��~�o1��2�R����n�8����bmn�C�Ԋ_����E��˳�GzY��%�G��+1�WB�/��[��bd%)�V�cBG���6`���c�rg�1�y5��o���0��XlxVHYEB    a19b    1f80����(A6����&�"�
]�-M�j��N�H���o/�9�O�ρv�y!�\���ؑ=MC4��q���8��D�_�Ζgz�f���%�������6�"�2S��=�Saw"c���� ���B���5�v(ǃ�8n��Q�$#݉r&�W@&{?��h�&��16�b%ʣ��Ö(�3x��*O$C9��Q*U�7�|�WP*�2g)(.��3��r\���] 1�6��J�
� X�Ar���0K���a7}$Z�L�H:~��d+[��W-7{1ML����Bl�*^?BF�~U9�("��n�u��=߅�`�.�Mm�xk&W	 �ʩ�Y]��}���P�|� xʈ�5�}q|�/
��p�e�ԑ�u�YT�y�0�N�#E�p��6�^�ㆴ�S�3r���ϲD��4T3[i�˭���s���<p#�b�����!�x��K�:�s������,\h�I��W7���U!�5G^���V�fnk�AXDM�5�����u3�u�}[e�vp&S�L%�E�>4*�o-LRW98�Ά밥�`��ر�p-&e���%���ڂ<'��t.U������@�Z���޳�L�Lz��-S�V )Z��h��9���.�Vxlkۣ�xH�v��o�mQ#E~�ߜ]H�1��lY� ��u�E����'��Tx�50�Ri�Y4n���O:6s���Z����?������=c�$Yc�QR�I���Ao�x��g%�5�L�<� ̇�a����CsqnG�&�,,���ٟ�D��}H��:B3]����Z��C�\���$���[����Ϝ�R/��R�W@z	Ķ�+LƲ�u�N7���jI���32,{h�Ҵ�?��+�����W�W��N���Iה�ۏ�A��	Ë�
�F-�I�*�p.^T��rh��z���,We�����L(2��(�b_8�PO��o�V�Vd����=��~#�l�J���6�N
Q/c5�4��}�'c�,�M ��(�dYvmr��ndb� �(�Õ����W�l!������QL %���\,y� �n���n?�-�d�pd�хzd��NC��z�9j#�mӄ����	?x��Q�����׈4Kc���Y��<ꋓ<(���7Xy�[(em�v�/��(Dw k�2Z|�����@��<�iڷe�BD4j-��k��c�� %��5���	�U���59�pXv/e��@ޫL$����Ϯ\u~�[�y�'Q�aE�0�G+F����.vqL*��m�\H�=g�1Z�����n���!E��#p{=33��ڰ�)'q��Ŷ�Rz���j��QV�chb	��<^_��l.�g���=�T������0���/
Nl"�a?��#��j�\��;bL!Ƥ���G�<�cUe1%*�w�3��x(Ƕc֨��?�Y��w=�%} #�F�cX�bub�
}q�"�49eQ�biʛ���x:�U�m��]��R��E
�[�LnĂ����x��
恍�8?�������#�(���hk��+2+���j�JKxa>�a4V����4����z	��9��q��!]��!�Uv���Sr��6$���o1{��?�X��@>���4�UGc��T�~6�x�3��y[�c���)2�O�h��ܐ3�Z���F���R��$]ؠ[��e!F��(����Q� �-J��d��ֶ�\WX��"y?$��!���Ѹ.UW��a	�pb�>/L�zW�܈i��E@��Bd�g�@��'��3<�-:~,%n�"����/a�>�5YT|a[?�"���{+�(�/i���\F�L��B�=ቩF`�S���͆���ȍ�ܫ��+�D� ���@�w{&k��O86��ך/ٿ�RP�+'l�C.��&����>#�~���fxP��>J�o��4s	k9��`j;�OҐ��ތP�ѳ]2�c�������U�"�|�ߒ�?ei�a���Z���g�T�w �M��@k͏�FE>��҈.�#e#}ܾ9��1��-0�����tDL�=����ߚ�gX-֋,$]�#2��UO
��2Ձ�jXF�}��x#W�x�t�,FHG�x��N��R�xX��K���
O@���J	:)�9O�4c�;fG~]0jݾ{��Cc���[U+�����Y��<[pjs�L�'��n��R�^go1��׬/T��¹�2�a��Ǯ'+lX�a���-��f��DtL� 5 !�`�P�4Ҋ�[Py�rva�$�U�gjol��y'zf5��CH&�C�^WoD���Q���F����pn/�|,�&�FQ�ά0���j��>XXC%�Y{k	A�,�9ǚn�).�6���l�~e>�ؾ1p 0��[$&��b �h���9h��N���$|##��=��Ӹ���*�H��.�r��C�SQ�IT��+9B�z�@���3��#��.�yU�
���S}Tm]H&L~(�cͤ�c|�9���J$3|8AM�bh�8[�2s���i-���%���`^�)%��+�������qZ�rL�Lo��b�ϱ3��QS18�C���UNs��&�bߋ���]Ǽ���qTW����z~bn-U��lj�+�z�Y&�O��-��*9�����g:�	��3��P��oisG�iN^�������v��yv `��~T̃}��.�tM�H�H�"��z@u�(�;N<�!��c�d\�����B�WM���&0��d����_��x�_��BN�i��j���厧2M{��^G�X��nٽ���R�y~}��3�k�@��!�B�� A��S@2|��ҥ��Ag}z
s\u�Ҫ�����8��^�k�em�m�9��6�@���,��@�b4j�=~&Z�P)�I�;��řI�S)��Q��u.|B��mQBWS����ӂw݈vl%�o�6����w�З��q�7�f� Q�H�������Z���Oʣ_9�_k)F�]����>Cz�ÂC��E1X\�W�iw*U_U�)B(�@��HnLXu*uJ<r[�+lG�����5��Y�ژ#�#Y\o��ۚl'ځYl��}�E. 6;�i�zR�Y��������}��b �ڐ�䕭�˸{P.�ة�Y�~��08}�!PS��T�p�l���?I����
`�8���|)��G�x���g����)�2�wVu��6Q��"��7:^SzwC��ݪ�R�Gb�	9RYJ���/Z�a�r��Xn����T�Y5�K���P�]N�c�&'�	�Y����?��"v�Jyk�/�@K��'��#"�;�Ҡ3$N�@{���R�þd���6�8ܮm�m�DO��s�M��E�ʇ����鎔��{_�hN"�'��ȃ�ؐS~��>q��(���$���μS�i���N|��i~���4/���'
� n�l�9Xe���Q9{��.��~��B}g)T�:iq���j4T��'��j>?Ǽ/�`}߭\u'$m@-�7ln��C�]��"���ĎJ,��Đ&�|�B"��\�m�m��/.x��V��AZ=�L���������Ǳ����,�[(a�i�e����>5�j��E	��V�}0Y~�����!y	owE�("N!�������
�L�����%{j���l��"l���3��?��KJ�M\}/"�xZ�>��\ޘXf
W5P��Z-ӳm�������1�#�1%+և4�DD8��*�K���Û@D�UpX�11�M������Q�+���0��7>�ϣ�`��)�A���p��<D8��=}:r�j��[�.�b���Lf?j7I;�۲��j�q(��9W�ks��yT��bة@	Ud�˵��
�gB���+W׏-����H.=��Ӗ�b$]�
D�3�)��v�)����j� 7����ɨA��)o���,�J�OX����A:p%�m�]x>�;�=�^gOW��vgpt�d��P/�i�3�m���4q��Q*x��,�V����s:�AB�Do��w�ֱ��d��-��Uw�?c��K���p�����wx���P�=��^L+�87���30��r ը���K���!9>��8I�Tj󃬻a���=�,�4�V<*Lt��6=���gu�y�NV��rpQ#���K�J�$N<c�}9{���j筎˖�o��$)�$�0�����z�n@�r�#|�E�r�l���/��M��<\N\�䳣� �[�q�%�������S� R���d(I��`�ZL,s��|&�)�k�v��Td@ �P�T+@W_D��"$��p;�oY��'to����'��\�1��d�NC�����2����ovc��C�%�C�W�P��$��z�v��d�P�-��Ќ�����\r�/���7�|��dB��?�҆k���ק~�ǘ?c�W&����G��
n�ÖX���s����v��,�7�v:�����`hH׋�9�ϟ�.���h�e���L����	\2j���?N�n��]��0 �\�+a�GӟD�)sr�m�W�Ir},�1�ö/������b����U���%js�����$��!>�uqZw��\9M�����dD���<���>W�K|���+\Y63Z�ז�˷���/�mf�Ŋ�r_v>Z�������Z�={�6U%Qn�邉
�E�y�����/�����._	R}>y�]L���k����dD��TJ�!k�k��о�)��[���E]`����0����Ah"���9�5��*K#Zڕ�5��&V���,��Ok���?P�3�&:��e�VL�R0�|�񗨿�iT��mDbS&]�Y���%��n���U�ْ��i_���Zz�iT����0.�.3o�s�9��*]Ү���4<-u�AӪ�á *��S�^Յ����[d^�j�L�غ�3*2W�E;(�,�b�+*;x�fD����0J���:t��3ʌp?�^��=���Տ��������о�͝����X��;ߞ�tRVC�_[?Hܴ|1���ىXb������?��̲*�،�P&kT�A��ͻ�ϱ�(l�-E�ܓ��kN�*�f��l�k��6��p�M�
fV<�F���F����ǎ&YKO-~��d��L,�߲`�<�އ��լ��@���)R��`�t�%��g�/��}QG���Ŝx��Q�GF����J)	D)�e�u�>�p�^�S_�\l>��;ŝ�֫�4`mC�˵	�\m�ԩi�3�̦ĵ�����Rh�����sAt�����.�rɣޛ�Fڈ
���|�'�D�$�7\�����t4�ȏ0:a`���G�v�H�������%����·1����3��%��U�B'W�|�-s�ĉL���B>{�Ş���.��^9�0�<��y���0��}@G 1G������l��+ε�i�����V�cQa�����!�粗E3��eؔ1��gy� �k��B�O?�����1*�5M�1�te)����x�f�[vF�V�H�������)�s���O'�Oݞ�6)nD��E�6�A>"��O�����8�2	zV��%�h�t*��H�ӻ�.��r�i�#�>�C�"r�hYH&8}_�Se���6QR5fN�_��hr�H�A�D�l�2+��lU��s��*3.�����U4�U��j�N�]�@��k��h�*-�cTR�g_(���rQw�p"� 	��ߦ�Ǣs��&�|�.�Rt[�+&�X�z�(ң�t��N��SD����
-��Pl���ް���|��ۿɨ�P;yo ���L���� ��l�Ur'|":(\�C�ý9�4/t#V�k���ﴋ��j�qBv�]���J<�&T' ? 9�_'ڛ�Ɋ&b�f���ky�4U1#�i$�^x��1�A�?�ge�)a=;�`�˔�%d*Ўh:C9�?���P�\4��E��Q�~���"<=!3�&�˻��7����N���>�w0XK��2�BWvD�C�Q�!#�D�� ��5� UK2�x��������۳����vP�'�^�)�m��g��I�+�]���jb�����T��s�0!�n܊���O�������4ȇ�y���AD ���v�U����CL��w>�WA��d�$$Y�9�x|b-���Q+ZA7�����n��=�z�C/v�:l��^��*��#.ٙ��A���Ĥ�d��0o�%��ǵ �R�y.uf��RG�C�"�F��F^e�<-�G�	0�}R ��~�`� V�B[�]��Ŝ�S!���T�k.*�u��X�����/�y�L��µ{x����ԓ�:�q����[�N�_�,��_��Ӡ�[���;�Q�i�\�A��f���� �0X΄L섚õPn�N0�6ց:!O�8u>�Y5�E5J YT���x���|'��f
O������Cq�"�/SgC�2�QUYC����ȶ�4R��}��za�d��8zN��3���G&ڏ��t������|E+:�����[��hk�*ͣ�I7�=�_~@�����è����B�x���)�w&��h	��;�^P�9T'�=]Z\ٔGS�0(FͽDQ������Tn�ao�f�Fz�S�0��䍥^�뢐�&�X�ah�� q"r�r��h�E������El��R��zC?s�l�x#���dYL�nt`º�]~�����C�kN�����\r�.�<^Yi��EE�<�\!160�!)�����ewO����$�K����w$z�񷈕��a�*
�2[	[���-�u�O��mԨ�K�>����%�>lF��j�"3۾>ѥ�AN�xg^���Z��s�v`E{J��%n%blo��8c��Xq��	
kx-sY�Bgw6�p���� �:���߭ݶm+�%�E�ؗ[�M�K�Q%��0��k�˶��ߑ�&�QrȨk¤N����q����Y!	�g�q�s˳l�>�O������+�p�~r7ޫ��yU���£\Hϙ�$y���2CV��R�M����M~ae�C�{�Y�Q�$;�Z�6v�n�	�f��8�R.Գ�H8;�'um�@_�{ۊU-��m
����	�/lJ��0����a0d���@,Ƞ�R���D#K=�e`	����ܚ}iF�����:/<E�ԂMp��|-ϓ�A���umږ_��qQ�����8p
�-\g��;G�Fc�Ȕ�S�UF�F�"Z��*Oy�6�MHVB&TE�L���h����dSb�t�H:�ʝyK1�]�d2��Ȫ��m:�������8��_h�9��u�K�� �_�7��XTtŮ�c#�~�M3�o��JFj �F1���kC���B�8��i�E��lֱ�SI�;�O� ��Rq+���b�(E:��ǀT�םK'xA�����%�yԦh<
^�1\���f�OCR2���ة[M��e�t���3\�#lk�AR9א��*�n���A���iU(k�����3#IX�)|�B�^�ټ%�vK��a�{���u��(z�KR�H��	s�x�x��$��}D�т#��BQN��yy�"4�����9�'�8U�r��\6`��f�a�˃�Z�����/���J8*��������3�5��$`��kTC|�P*�o�\i9&zs�H��G7����x(*A�Z�h-� ��q�n�1����<���Ǔ}������w�3�R�����V�#��O��w�%�u�}��@{��q��o3�
)�7�!3vJ֛��C�B�Ҝ��pŮ/
�����G�h�v��L̶&�N����κުV	x�qS�a.>��ጸ�!J���%����E�D%i�B���z�ǟ�n�̛��]NF�l���՘���q�@$�4�L,�	B-���B�a8O9���^\o�:�z�57F�_|��Y��<��&jQ	�6u�\+1_��VJY��H�|_<�;֘���pZk0"�$S�J�%l^k��I�/�K�g���,���Oa/�4�	'>8qj����I�\9O�ٽ�B?�����ָ����	� p]@B��] m:��|