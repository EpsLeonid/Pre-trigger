XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���?�/*������mD� ��kE�¨��H$�k��6�;º���e��8��q�b���s�p��;�k'3�� ����=2�pe$�=r,ŇXW���	Ozb-��(����z�� �3�F%��S���M�[ n��˟�8���}iIcs���H]��]:u��?zѾ:q��z�w;gƉ�4�L��ٻP	�R�&�R����L�?�%�C�ڣm�eaP<��T����]�Gg~`c'm������i���dU�&��?�>���������5�E�˻�ƈ��H�ݡ<�%-2
�-�	�x��ޜ�ĄF�]@(��%��DW��"+"�D3}�[؁��x�?6��E-���G�5���D��
�ݣ��Y+��౪���?�T��O��i���}�8�Gɪ+��l:�+�7��7�!_���W���6�SiR���kO��gy�i���ݑ
�@7N�����ݪ�g_�B�qd�^,ZH14|,
�L��q(�g-��Dxw��~=�!vc��C�Wܢ᧬+��.~z�V5C鎍(�!U�'���kw/7t�pg��]��J��?�I-����g_�_�?���U>���"d��ZN,=��|���="���:��"�l���Aӊs��i��x��\�VSE}^o��T�OЮ�����R�_�����=1�K ����#T��jL��KJ����I%��(R�2t0B���HFH���n,G;O�WyVi��n�� �H�?N�����L������XlxVHYEB    2327     a90���+�.ѡAO����s��b$��%@KK`�N�k���n�(	Tv����F�<F?�?�d�y���)�u�,9I��[,���:`:��Wu�	l��"�FW9�:��iTc��{��I�f�v}N���tt��,v-�ݔ�b��{݉b�k���{��#�#�n��m8�[*p6~�ذ���V�~ԟ�Mq��l�����'�\�)K�GU�p�P*��[������Tb����Ld�s�_n������i]rZf�;���Yt�l(W�S�m7�NФ�*���XN�g�k�޻��?������s��y�^AL�g/e��BC�����hh���d�iN�!�jw�5���;��Ew�Q3?������1�JAqy�/jv۰�e�ެ���X-�F�������y;W*XZ�,02�F��G�,�p���ѓs[Z�v��zV�^R�+i�Z	h '��^�-���C�+��Y�d��j!����"�'�����vA�c%�$h?��O�L�^v=�Ċ�y㇛~�N!M��L��xW <VO{*�I��=DX!~2\�r�21�Y�ZMc�E%z9S�=��Τ񒭙��Nc�
Y�m�YH5q���Fy����v(�D��TK�(u1�2^�fMs.�I�wn��Eg�bW�I�W��5���*fb4 b	�r¾��òׁ�Rг�{!�]oE[�I��p�#"̃Q�����q��	=^��҇]�sB�#.=� �l^۰��삞2˛H�ު�� H�S9>F����w�����Sz�`ظm��nE��=f��0��a=.�K/��0i��ф�\�O6'��8;+�b��R�E�EFT��%�`��,���
�?��1L/N�4b�<��Yj6p��h�hL}k���,0��^�:g(酻�I#c�z���K�9r�o�u�J�L����l�ω��ħ��.�9�V�i[݊�G��˟A���f�]����r�v��7�:hw\M@�Ǿߖg�M��'�p'GW������a4 �w��8�i�`�xw%��)�����9�y���7̵�{R��Z��p���VCpFDj�~2A8�}L�e�-�iUXPO!i^��G��Z%�?���dJ�,^��F+d�Bll�m�ئ V�k�|G����!���Q�<�;�%��o�����ŀ�$�o���
&:������Ϡ�)�Ë^�S�C��z<⃟ϯx�!�3��l�,�����G	�m�~��������er���E��1�it��'3ߓҩ}�\$�䦪�t	ƶSȘ��ߍWMN� �voc�s9��;�J�bo�ua�?l\�~a;	ERz�2U=�)PW�i��ZT���s�!˹U`���Y?�L2�B���Ă�'��,9_�*�;=怇��)����ُR^Y�=c�5�}���9|¹w��Ռc��6��蟬a!RG�o^[V`]4x^S~�w=2��0�������R����~�~��S5�5���.H�=���`a\���s���u�6K=���`b{�����ua|����Ia���C¸gL0.���F��&��7�{aV�!�$� ��Szo)���od��P�'(�n�	�V�H�f� �8a�Z{����*� z��Q���
'������F���-�pʱl����k}_���}���cJS6<#�S)�gK@T.�]f�x4K�$�Q� �{�;͖ܙ 1�oݐ+���Ͱ��y����~�ww�~��X��3��Ìf�պ+��^��.JՏ>�r�0�ݫzPeܘ�l+�dB�Z7:�\U�uZEH8YT���EI�N	Ȁ�}�!����;�^�#�sU�����֗+Of���&�&u
ǲ9�x��<�P*RfZ��p�\���_g&�d37�4^����\�J�|��7���6��R颛A��ң���3�TTc�b51?�w������1�4��c����T���{��K"�8�[G�"�CC� �'��G�<�8W���"9�(�H���[Ii-�ģ�#~�4�kQI���;v� 8l�\���cȽ4���?_�H��G.����d��mAs�>8U�R�H��Ed>3pZ�����T+Տ>}a�{�eR�Oب/�o�há�t)0 ��!vSz���A�a|NHS���1�lm���);�����]����B*���tȠHfUPKyH_��.a�W����	��<��OSgX�@��S�ވv��,j_�h���c2N��V�Wt��(m@�N_L��޾,�8Eo��Pt��^"���Cn�D9
o Bαc)��Ӧ�><�h����8Xz�+kz����+�����c���{��!_TZճ�>N��͗���lk(.`�@��8.��$�qM�w�����o�8׊�w�!�Ճ���~���s{C��x�(���V����P δ��$ƫ��Y�o�
�[�s�֊)gȎDa��I�E@���I%qd�ܙ��xQ�Q ®�0�zghyv��}����ɓ�E�Ь�]o� �yz��-uE�zUnN�؂��(X�����y��O�B����=x�����S�I�P%A��ߢ�go�L��?�P��G��88�ގ٫���KC�<��b��K�E��O���@�M�ak	@�噤�R͏t���Zz4�k45�k����xZ�qkbq�I9b�
rk]u����4�݈Ȫ���l