XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� �-HxFŪ��izM�k�P�oD��ń�;F�y�oG������X���U�g�x���L�èG�iL���褶Y�%f���I�<�p����~�W�]����@�	d�5��}Z�9�U=-�#���/n��/r#s�����Ѻt�H��HP�e���a�u�N���2P�#tV�̝"T��C�UT��v�\t��0��:�)sqI�B�g�/��^�5s�����v�jë-M��=unػ�-�'id���W�h�����7#��-`�T� �xOY*�-�/
�t�r�Lh��l��@��T�8���7z�=����\v! �E,�A�/Τ�VQ:,#�پ�2�e�+��PD���9�yi���YoX�AHYO�gR������8�j� ,���T[�%#�$�|Z���؆���e��x��$��$���%;L}��n}C�$�E��{"(p�Y�F5��Q* ��T��������iwԛ��|@.���b7�����{���c�ޅ����V*�����FM_D9�� ����#�$������F(+}��d����kP����A�����w��[����'�?Y���$*���wڌk�f��;&~M��V� �f�8"E(�P5ԗkYS��:�`���?k�?�����:�9(���O�~	�S''��x�OSH�lk�O$�~"R�e�2�M��*wmg�1&���TsW�]0�jF���$� ľX�1|�S�8��_��,�y��Aȃ�(#�|���4�XlxVHYEB    7a7e    1af0��Ŋ�n�������֏i����x�3w8�.,TPe2<���q�XS�	/�?Pe�@���KAq����Bt��IaAn��th}^��ӑC��>����霚\3Պ;`�a�@Dt�*�z�L��p�t��I!λ2�I����E[G��Q�.I��/!�?/�h��	�8�����@�P��9Fޔ��b�-�Ҕw���t��'	!���'���?Ď����9((9��-�^����~������V� �RH����w�{�xɃ�3Ã���y����u�[�B�4p�_������9��?�Μb����GOM�$�,:��ۋU��"7��PV!Lu�R��)����Fn����� ͱ�L�A.F�,M'Y$̋i��|�̃�ޝV�T�x�]`S���r�Y����p|�ʨ�
 R;f����`Y�s@�q>`���a�p�T�q����]����Kұ]4x���[�"�����"F������'�$J�x���0�_�9sVCjزɩwˮ}����K����Fay�����[�Ǘ�^��e.6�'�^���#
O-h?mMWOW�|�:�B�^椚�N��#g�����P��ZNb|x�]vb�F	�%�ʝ���g�ҳ���g��"ه �̏d;o�eh� ��m��w�tX���	M�$F*>n�Cs�^��+�>�k�N�3)����I���J�Wq`�$ �ÖF���`��s�@�A���,�У�Gנ�a�<�`��#��d\��֍%���.��8�ư��o`.<D����~�Fj�3��d��������n���9��4�B��������^!17�/�r�HKj�ngGܢt� l1���Ml�O`˞�?XZ�(u��B�iZ� �м�$���W��.�رɆ����A?�L�Tjh-g�  ��5Lp��z�m�g�F�y4g3!��7��[�*`&!�U[E;Ph���6��#IW9J�52�J��j�P������� �C 񗄐� �������z<ҩ�����J_K�H�Z�ɀ�x�H2=����<xEgo��7KH~io{�C�@��X���2�a�ҏ?�vv3��93�&���fd=,ݧ�o��Pa��Oj�x
�H��<ԯ�Հ���H�{�G2k�$�i텠y�62X�0mkG���P����٥F>������7�����S�e��@�� �N�T��\8�"�9҇'���{:�s��@%�-$ָ���i-\�-��&}K�>�\LM�\�(a���9וNd�E0	ht)��BrQʀ}�W2\��r/¹{�/z'�!�!L���8�ܩ,`�U�3�^��}�c_\FJ�R�1�MN{�B�����p���ʣ:uIt
��NL���R��DU�A���M�"<���J�$��F
`��k�hS������9ě������O�Ϡ����&�����SĒ*��hU5�e ��7�Z�M+���ff`Y�~hY�陘��n����7�r<�C�25O�$�|bX�W[ݖ�#�^uh���aU�c�g�?/k�V��-< ��`�ō��L
�.�ҍ�+N@;h�u�c�	�׷-�>�A��tV��Gm����N�D Q�W:ކ?�h�d{Q�8.��p����3U�6.���|4JEG�F:+�����b�ҟ-D���TIG��1~:YZ�C_�Jjͳ����v�}�v��n+�Y��ѵ�b�k�^�ƉF%��N�T�g��آ�5G��ۊD�y���O�w��*	(2B5��c��xJy��|U���Ζ.E�Q�[���1��@���%�Y��b�e?<#g⅁��p�"��wT-(`:u!y+`_9�#e�/��V��;a#";3�u�A� �	˻�c7�'��'�p�~un�e�&�[e�E��tkr;�׾kOG`9;���4p(p���r���!6��(�F����F���G^�c�w�Y��v��2X��V�a�2"�GJU!?$V�x��J�k#^�-ud�7�zq���;g��5S��&n['���0fǸ��O9'7�1M�i�g�5�����i.��ϝ���+O��5~0n���$G0VPw_���wV�-�$���c��G�m�fS�*�ͷ����N�9��N��Y����)�\�q����� 񗲦�9)�=���<m�p���J�����F�W�6��[�N��}������i��Fޱ���V1p��3 i(O�Pc�_	��G{8���'8�~I��a>[F�I[�3ҝ�/���+���B){j����l�[e��w����U5�������<��
۹;�cs�반�k`@t����K�L(8�/��πܲo�?괵o��^���8��wu��~nW��g|�Ap�j��X陵!@ �מ���J��F�£K��8��kf�\0w���;��Q@I-" f((��P���#jXʈ\���Q������1Ya;����}@����;�ҕ̵"{��,�SC�ނ{=R�G�-`�D�%N;��:Р�Wc5�R�@�h�
;�!��i�!O�x�V0s����dm�� HMU'�6l>6:��:b���x�L /y�5�+4���ɩ+�����'�;hi65wgF,A�o�@��a"��n;�|W�ў��,�ۂxY�1O���m�-Z��g@̬59V�@��-+�î�0��К��m�ϞZf		��}s�$��v���)��ģZ�G�i�Gɴ�*���?v_�
gW!�QVk���r�D����_]`�W�(�E���Y3�|ڬ��հ�=elz�v���HI�{M����U�y��Ð�l���K��˨w�&�&��/-��;�CL�vգ��c*��IR�Ͳ����yj�+)���t�&�`2Q������L��8���p��LXV�Y�n*���m���追�n�`:^ov<2Q��NxCf*HCB�}����!�D�ncHo
T�� ͱ�z!�fq�����ݥ�)W�#z�}�M�r��rJ�=8�!�4�*L�F�gt���ʃ3�T������."��GƆ4���#(����HU���#��.:�ػ�u�b�U�E�N	���+�ˋig���^ݠ�����?t�v�P�?׾�Ʋ엲�\!).b��-E�$W֒\�3�[S�6=c�4V�����G|�BC�i&�A�u�S.5�&_I�ڀ��Ֆ}�am:�,8k�t=d3����:q�r�o~�k�l�0$���$��P[����P��2e��4�Sfn��>u��|n�!���nm���A���HY�
�&�Yi�K�lߵ*�� �F�XM@���Pg���T�|��R����j�A	�f�*���PΉ�%Čь~�A0��B�3�O$�L��ߨ� ��]�1��P���'��C�Fg�n��d+%p���8���S��[�_29�Ԇ�*��W4��J[@�1iM�U�����t��C�!�����|n�s�������\ٯ-5 NH23#s&wE����yEwp/�٤4�-���#6e����]�2��Q������+�T$�2\25��-k�0Q�밫Tkr)�-3e�j�u�_ÊU2�Te�n
Lyi.f�2�����Z�O��O�Ht�S���0���A�4��Hmp+�H �Y��8��K@3�#��X�Jڔ4���D��������r�8�d�p���s�F�̒$���o�?nw���W�� ��Me��n�6Mo�A?�oMxS	GL+:�O�<�=�4��s}�Ss���I ?途�d;�ă��׸��0�)�
6��۝\]#4��1�G���d����}���8ZJ�
Q%W� ��:���c�m@ �ni
��9u���h"���9���4��_���Ԅ&�����$u���R�O���eh�&R��1�m� �=�1tA�Vna!T7xOg�b������{��,�>�md��J>)��� �AY��Tt� �+��}�{����� �|����ѝW�4]�ɇ(��*=�Tt��@�6�ă�Д��
����Z@�3X��鿈AZKG!U�%����5�g9��?}11�z�W?�Nv�ʋ�ݧ� �s^��y�Ҝ�hC�x��X@�j�#o�E #�rl�C_;���s�-a#�qi��ob��A����")o��#�m��Uj7h�V�����苒�1����2/�|Lf2���cC�4=�{g���J{�|�JR�9�T�t�.��c1/9�?�2��T�"��Fֵ�3��Y%P��*9dS�}D\�@�b6�W�+���_[��!6q���:#��i��ڝr'u�J���d�n%�S/U��cs�!�DH�2Ң$�=��7sB<@��o�=n�k�ԟz�4��ঽ��kmq��=OlDtFW
��� %d��d\,�����L�]�.��b�;�ʹ*��R���圯%�i��e�(U
��}S�����C����*�UD6P�ʪ��f[��gW� ΢�Ē�;�>��|��lk�m}�Yu�J1Fc��jx'��o��\�k�����o�۶�n�k�y*�z*¯��ӹ����aZ�4Pc��,�|5�AE����6(�5cV��`-T��cz�G�%���/�Z�/R��ܼ~���,�S��$��G&h����ԕ�}ʑ����%�M�ak�{�:����tUM��{c��(e����}�)#ʸ�ԣ��oB�䩠KU����,%[�\���7�T-�K�.g&H���t|.���XFi�4���r<Vmx�I��� >���/P���@iJ��G�-��m|'Z�Վ���y�ʔe�D��?%S����+��홙*���>oJ)�������9���uH'ӝC9�x�)�)F5ϣыq�ɞ���wV9�o�@�P���l�F�q��BA*�-�Be��p���<�gٌw����
Aoa�պ��bl�l!�,��&Cq�µ8�O�'��zF���Ej��P��h�z.��ظԲ�%LQ�T#7�8j`ѾE�{d���E��Q'5��:K�t��PMrA�#���@��V�X�h�p)��SA*���N��L�e'����W�>�'�9����BkX�zR��#�C����Қ^�)��u���N�v\��AE�W�"���A{�����E|ׁ8�e'�>��K2f��P�C 2�;\cOL�װ~���ջc*(	t/���5��)I������c��Ŝ��\cc�}�ے1�Ȇ�cۙE��2@�9 W^��=��24KT�%sT�]|6�+�0]LϪ ��� ��F�"w��®4F��A@{���\��=�F�[p>�r�C���M��4+eMpU�-K&@bL���X�\+W��g�IR���l������@O�Sq�x>����(O:u��VF>݀�?⮐���NkC�G�\X^�P��C%T�2(��%{ǯ�`,��xo�|�V6�[�SJ�kSS�R�,�N~��+�烳vA��Q�k�������7�"��Y��t�Su2�fu#IA����@_�#�Sx��(�*t�_;�U�Uv�IXևn��U�D=��+jS��Ps��5���$�g������)t,)�W�yx[C1�O�x���e%��<�
{a��m�A�)Dt��۽9�4��cD��ek�s�VFC'Z��sV�$_׼٢��8
V�M�6?������2���֝�R�?]�����m�u��?�FP�IuW���6XD�xP�c��|�Д��݋%�"Z?�J���7vPH�u%��
��1��(5:��B	����j�/ַ��K P�]@+�3iO��S|������ʃ��tK? ��I������/���h��π�ng��N��^�Ϸ�8l��� ��mŧn�\�3i��+V�
vc��h�C�m��pTāq٪���J�y��N���*�D�g�TmG�l���w��2#�|��חZ�an����D�1���W�BJ�S�ڵ�8ղ8=��"�j��y�!;l��uK��J�+[2�1e���Az���Y芊�U���P>�%�:#|�ʿoi�VG
��d`n�ʈ�
�%h�-�,�pA!Q�`?z~R������xz�C�y��k�Y;��5��6p<�y�Ŭ�ѩ�8��k�;�>U5��:�)&kL��<�7����hS �j�7����(m�m>��Z^���}�2Y�#�=���h��K`=��S_���3�i.6�L�
�o�\7�IkK[�
����=�,��o����}��C5)�_��p	�B�y+�*���\�Ism-��7�Χ��=�D%-[��	�Dm��N�ǥtL3�m�=1C����i���g��h���X�=���gaثky�1{.V��6�����=��o1X�j�0�$b� J\�w�v{�j6��[�&���j�]�S���o]��L�RMs/���[-�FZ�ӍE�c}e*8p�.cO��D+F��B�Cvz:��s��~,�v��7�>}q����u��	[�p�<&8~�x`����j#�)��F�G0�#�����ُ�z�d�)��b/�����7s�
�{��{!.p��O/ت�^�ej�����J*vz��Pc2��b���G;sqi1w �Z�$Ӳĳ=���{�c�a<���}$��"./����{�=��<��gJ����}��?�c����2��B�=�ɪ�I�x�B��9 ;�]�a e�H'cj"�xBbP�~���<���h�<�K���9�b�~in�h����uK�O%��9�Ul2ր�Hx��_n��x�;�\��3v*ŭw��Bf����*h�av7C�	J��
88-�_�_�\W[v��1o�G��+}ƒ���d2�