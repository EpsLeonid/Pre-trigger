XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���]�~�Щ���o����TL��H�����W2`ٓ:k���_Jа�il`��hch��Й��y���b�YC���NCW����S���F#*;>[���KaS����1�N�rJ���y�&�|�!��r+�h#����i1�b1en���?�������xP��,�}�����u��~��gc!C�ѦapN��}�ǩ�qpD���u���Ts��N��]���C��3��,[����+%{I�BL�j���,1ܩ����C!z��g�Ĝ.�fS޸�nʋ7!�~��#�8�Э[f�	Y�IĲiӹm�씷z��6�?,a9=��Z?�'"-p>��5�� �m��R�^O�@7С+���:y�2L	�)�{����qr%ĴO�B�kܐ���֟���񔬸
���,�o�|�ΡI�C<�vy¨_�.��72E)%_�5�
���#g&��>���W���L�+�^ƈ���~�2����
ՠK}AC���)��FV���~\&�n�����&���fi����m�0��0�q���ZH�K���qM(�S+\��|&������4B�J6�ߨ�O�� 3s�)|MQ����(�|��n� J��!��w*���Y]����c��,zDм^@��x��Nf8]TM����S�z�fh����HW������]+ڞ�ܔt@]Yv1�����9}�$4���a�s�n��:ʹ�=hƚT|1\��D��pҀ@9�YXlxVHYEB    2442     ab0���D�ڪ�O�Z��5�0}�7/#���.y���Ů���ɱ�(��hZM��1
��x�!4O��?���py�z��UO@E��	��ㅿb~��WS��"b!����a��g@�����/��!,��,�3/����2�N��L�(�s�V,�F�\)�z��� �
U�����,����U<�Qy���S: �h�F��]4�cf��l6N�1�9���\�&�^��ɆU��%c��M�F		v$���U�g���n�HT��cT(�(�j�R0 (	��	�	�Ԣ7��P�����I�6��l����$��ԏ����Z���V�[>Fw���Z�Q>�rA���[��7��r�f��q��c�M��wПD�ϏP>��>�n$0�Dx�+����80�m�������-w�"X��u#6��>h#z��H�<k1�)5�3�τ�~�yr+C���+ٖ%pu1�7�6�5{�3`C��8�� ��V�k�<U�WH5);u-��z���îh�5���f�Z[̜ˬb,���ã3�CtIц]�q;��⪽���/������f����w{�3*8��NJ��'�����4u��i�ۀ�w���-=�1�!��]�z��c�٣�*�NCu�+	�\��I�����,'�E�a�
�B0�^i�$x�E� ���4b>=U�8�H�92�ك�V�����۸�we�L���@~�7�, ylj��q��S�R�v_��Q�m7̽��E�?
K\��k�\&�MZ/Ov���z��D�me�z�3bjH`*���ݿ�j�<�U��9.�R������h}�O����O�f��v��V,*9��,�M׸|��֐�g�ps�| �)��7Tb��f���	��R�.52n�⺯4V2O�%+Hw��
a �%|��3º��%��S����9�����4��]@�Q��E:Z�y�&����,�g�$���v���@���[�:�D�f*N����秢�@�ά�x��3�����7u���Vdף'�
�FMJ�DϤW��U������;|i��.�U͇I��i�1����$V�XB
�߃{-�[�{>�B曢�v�7f�����/|�+�|���i�3ź��B�
�6x[�c�"��ܽq�ۑ|�SU�#U6>.�S[d�{�4�认���.�D������w��	D��?��h,We�U���fe����}�n%ԣ|;sڐ+r�,&�n[.w�H���_�X{i��[��!��Z�q��y`}39F�c�3t���ޡ���0Zk��]�|�ݛD����7�/�o��r��}���J�1:�Z�)���p�> 9�9��)F���s����j�i�E�.�̵��Ոg�UxK�R�f^�Ŋ�ȑL�W��S��~� �q(��	�(�k�#�0�
u��sb�=�����ɩȟ3�Z�����%Wϛ^����%�5Շ���T:�D"��o^r�r�� O��r�?�^{�A��EPS�dI�t)���L���4!S���),B�і���&,�荛��)iq�1�ȍx�H#����]TL~\ԦqE{Y�!@�R�E�e��H�%D�Ա�t���_��\�?:��ZP�~5y�#��&���Ž�ڮ�\4ǚ!��y�"�5̮4V�Q��_\�'A|'�L��֬�#�>�����+���,U4I����%�P eD�|���'�
����%��,�p8����#Aδ��i��A�i�N͸V���@�~Z�Zj�uX���o�Z��7rL�z�
�K_p�%m����Ĭꌀ ���~0����sU���xV#���Ս���oH�~E����H��t�w��u��䭮_���~'�cxuV畚�#�yؕ�ui*8�*(\Mq�������m6c�mj��t�$�(���f�-3��iϼ��7�;��]>�.T5�+X�ַ~��ƈ%y���ւ�,������z�4�>�!�t:��dK�Ww���zE@:Uhɺp���nnbIgL�(,djBD�Nun�����"g�^�H�=��-f����S��ms�c��C6y*]_����Z�p�h%Wa5x�ٞ��-��6?���&�0��>����A�����@L[�w>�QI\�����T��O@�mpA͉��H�{��ot��S���Z����YU�����������~�(���Z�(Y���(��L��?r��؝���6L�Is�P�:�W՞�;4���J��3e��#m���#H��9���!NZ��p#��撲+��|�G��Is�ѡ�&))^���D�~�!��U����w_�)�iϻK�Y)87��"�v�l#���ӷS�o���"(�9ރ�zOx��'�g��3όB�n N6��w.ڮ��<�ݵF3*H����%��ہ��&�������0Z�����\g�j��6�C���'�/��4O%-%���A�gb�d�M#��5��Qe˴�6Ͷ��x�v��~�aj�؄���HCP.����*�T}�����c�*�.V�2ڭ�S2P����*#̮�zS��zÍ*~�����o^[d�I�e�1qCLxBM^Fk��QΕ	b��$�1d�;�H�R�Z��#�Sw,��@;��7j̚���ԩ�Q���X�������̭��!��D�>a���$�9>�x�9Y��ו+���PЫXt���8����Hyh�Ń�KL�n-���B�j�?XN}t�k���