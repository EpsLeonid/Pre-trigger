XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��wp���c�{�R6���Dl����2>U��=��k��A�x��:��W�1�@|X�~T�$5xy��BgN�7��e�g,,Z�
nh5���#�;�7b�������9�]�uo9�`/	��'۳X�ȟ���C�/�>�.�����WQ����cyfAѩ'�N#\��`�����8�լ��8�ȗ�3P4V�*��R죜�V3H�w�̗�6e�~�vЧn�!���C��k�x�����#���:]�։��m$�vb(o;�!t��M�g�,�%�_s��0��ᮒ�gUS�XA�7��&���c�vBqY,�ezL��/_���NK�����,�0�{���_������Iq��%2�T!?J\r��< [���Qb��"�i�O�cֱV�7�͔�j �E��2�G���\�j�G��R�[�dщ���6F�k�(P��
*.����q�dZb�����h�R,�.��`��g�h18��ci"v�=�I?�!�N�k�X��ɣo�U���~[�1h�z�����]���J���9W���(�����n*������N��[}	��-�>���d[�7��b��ga��'L���M�h�V��Č��Oն��o)T|k�~�|��>� p���TJ6����7���n5���e)���*6!�Hav�S���,[����uFj:���eP3D?��Q�B�%)3�Z�-\�z0Ο��b5 8��\z�X<���@Y� �"��1��&�pT�w;f\	,�,��A.���a�'���&gT�+�8XlxVHYEB    3e0e    1150���v!KR��E������μ��Q���0�"���@���ߵ(�EQܨ�� ��#��B<1����#�y���U�P�Z��J05�F�&2n���p�͔1���'��q��C�&~�5���E��D�!�ڴ_o�u(	�����bMlD���5�f���<D�e��QJx����V���sWH��s�� ,}l���{�057�N�b=�4��`г7HN�l�
�w�k+��V��F2�L������ag�8�(�!L�*�ǔw~����P|(]��_�в�q	|}�X:���?2|�cM������'ņ�9.�����;��y����ȳLx
^dU���)]n�z�2�N�gπǡx�7X-���r*s�F�)�݉|�~<�|��qF�`����!��SZ��T]����gHŘK_�^��ȹ'MT3ɶ�𡯘pK�J���ۦ��}�k��Ms�Wi�:��6�,{R��*$����a1(�u�/�r:j�B��B�%�qGQJ���x��d"�����]�?EWR�V�Nle�K��"��!�h��p���E�ӚJlc�����"�?����xU�.��i�f�`$���U�����g-�{{� �� �����N�m\L@�`�
��&$�٘�i�=~Đ��>�|�yD7��N�Y�-C|�_sF>"~1�q
g�[��fh��N�S6���} 6Q��K��OfMF�T����[q�Ha�qp9�0\��b��֛��z�f��b{Yc�8c�W�����[�<� C�;T��fItt�+9���Ԑ�'vS��c��|AN����(�C�B��b�c��jb��ȿ ��-�#�r z��ݟo�vK`[A-�ړ����-a���6�ʚ�^�50�<ך��]IL�IC�ȫQ��}w��@�G:��� ~�q�И>�SFq�8Mo����C@�F��vj/���!�d'��	���7�I���v�=�@w�^�{��E8ӹwE����
qa׼�P$��)a�6p�����ʮ���I���UW�CDc��z�5��p��v�[ӹfk��k_đ���Is;8O�-��Vd���i(Aռ��,\ �d>����+��b6�>7����}Q,�ja�M6�V�� ��걙�ʒ��ڮ�h�������a����_�iԓ���FW���=b|K�ڡ�s�b{�i#�n'3�"�Rk� YK�@��һ-s���|�ZNd�b�t�*�s����a���JN=��� >�To�︽wv7��c^M,�����~�4�/ُ��4Q�OT����3�m
$8�Q'h��d��i+�C�t|1����[İ���WX@Q��A\�uJ&�ǝ�cP�o0�����=6M�����_���B��`y���$�)Y���x��H+��t&R���t="l�۹��H��Tq��^�䴱���5���Ȇ�r�W�B��RN{��>��
I���0�����r����Y(N>/�Q���?E�C$}�| �$��[ h�u�W�n��#�86)�x�:��J��4��$o��$�K����dL�:���4!}�'쳅FC}.�.�E����S0d����*7d�V�t�%�pչ����}L]��s�,�u��0��G{)�/��\+bu.4�!�mM'�:����xKuF i"���_����6�W��8r�p]� =��"'���I�e�]���_��htwW�H��L�F��&wJ�t��M�>��E�y�(�o'���9����)��Sm��ѽ�!����T[��T���S!����{��>�܁x;��w���k�D�9��os��BhqV�Y]�7j������m�
��LW[պ�R��=��Kj4mN��.��cw���|�&�`K��5;���|]�	H�Ű�;?J�N��r���&c���5��z�w7��a_�g�Im(7�9�M��!G�G��~�����؄zp*���'s�S�֌������LK��ҧժ`N��	�F� k}q+��G-_O<�(Fz~F��5 \i~_8����zU8��)P������~���}'�{{^���0�������)�cU����Q��J	�
����I��~{y����y�U6R;�(�]���<1CG,V�o Zثr�<߁�e@h�zfu]G��``q�g}Yb�A�~!`73�4n8���{U�Z�)�, �6�j����T<#6�(��w�z�X���
�B���Xv&���C��g5�8���O�˿QX���XU�iS5*O���-W�����@��r/�sE+z���dx��(�̮oA�Ȅq����C#�rW��ܶ�}Q^w۬���K`��AK�!����sh�G�=
AI���l�l.�{�*}F�4�

̦����� ����e_� 1��Y,QB�Mzܡ�,Չ�i,��^�Dv��x���<#�?[�16r��^���*N���:�T	3��Tg�c�u���T�(�˳$f�>bmfvT�����)A�%v��"�U��A��Tk8n�F�1����V�	8��Iʋ3�D��:G	��Y�H���J���E��G�ۀ^]�[<LD�AW��>�/`ad��E����""�~�*4��N��q���9\8���.6W��?�ᄍ�"<W������d8��ٵ��R�����ft����z�x�
;��D�Sh��M�3�J��u�c(�P�q�C?�rC%�<r�2��*�P�ΒF1{~��Zt��Њ�>��n���v����s�| 2��xLP�j�wl�q9��]
a�)���Q���;i��_�M�X�`d�e�$�+"m��v���.ہ��;Ģ�.����BLsaN��H	dX�q�͸(M����f�@�X�}�V��^�a�)���e��u�Z���k�����c�u?~?[�h��k��n�#Z]��2h)�*Ρ�_R����]��s��&�^TS��?�-�S̞�E���F��3����3WHK ެ����| J���\7b_��<Bd
I�l��G�A��=����!�8Gԟ�X�6�ɁC�쎄�Q�;�V��U?��)5�C��\ ��۶'k�W��k��)n��%K�B>�s0;��AW��s�Y	�kY���Clu8Ĝ�4��Џ�a*lP���;�Žx�v)�ob4+&6��3��-�*H��::u�������'	$E��)��k��2ތʄ��}�8����{
���2�K�Nמ����䫋E1��!�bɃ:�Rb�-J��*�i��9�X)M�H8\|���ax�����BO����9��y�땡P�J�]	(�YbB�K����薳�p��
�D�ANkX)<'W�w�u�J~P�P��ph�8�Kp�9�K��
���M\��3{� �A��k���%m:O��za�v%�l�!�Ȋ���@KZ`� ������/�wg�������A�i߰���^7��EM��7�ѐy��X�̓3SG,��i�OM����Y��9�mb����6@��O��?�f�	�<v���̋/��7v�Z��K�}�'1�>;篌��<i;c�Ù�Dr�)�����͕7T^�{A�|�P����n89�J�El/&�:!�bO߻�8�)�1�_0�O[�J:����}v��U�fMXZZ���L2렃>]���d�K�=� ؇�0/��oG���Q��ÒxiRx��e_{Eʐ�K���H{>c`D*���F3Ǆ�ώk���]�e�*�w� 2j�r9�<r���6�qT��tf��W�B\�
��՝L��}���	)��#�>�������	��KI<<��Ui��/7fw���E_�_������x�nltxh�&�A?#�����9lݠ�}Q�{��(�Q	�a'Օ�ᢚ�@��ʍ�����v̂�V�b����|����9.a5��?_3K�Jx���J��� ���b��Z�Kx��&=W�.���0�,	U�Q�����a</�m���چ�(4�)��WPy+L�ݤ<��O�1\��s�ي�T�Tc��5�4;�,��g� i>q���4�RUK�L�M�U��e�q�D7yQ~�Pu��Ƭ*?�>HY�6�ؘ��WܐI��M��>:X"ϚǦ()�'��)A�1݆��4�����1׹N�{}lˑ]�gp%��~�W�S�0J�yj�cU��Co\�JKB�Cf��e{K�w�яT�6O�D�(��s��{�/��<R�D�����*��i�*rW>0��θ�]Ɯ��ǅή6̩3���C}��]hW�{��\�X�r�ȑ.r6�҄{���щ@�/�gWhqN�pC�ʎJ���u9��{�T�u��+�'�����C������ZL�w+�~Ru�2,�+q����ۺ��g