XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^6Z�[mCR1��� �?v�fZ"�����u�s�k_{�*n�\�����si���Fc�/�ߔ���.���� ��*�I��#[�ja�I�� L�ɬ XĈ������m�����D�\ɶ}��~��)/6O����E���?�^��>k����;�����h��e6T�V�t����E�!�h�^������*�<���p6P��w����)�
�3���ó���
ٜg�,{h�ɻ�=Vo@����V ��	b�/l��k10	��u�c��O�6�N���p*]oP�6�:}���W	f]����͜���MYɷƌ��7|�-Yh��*y�Z��%P,Ue�}I~!�AK;���wC?$Ci�y	j���m�'-V��k���U�՟�۝����?�t�|�4��K�V+Z�TU��a���ꏆ����yv7���(L������4Du�<�
A� �.�>���%���7K�{�� �h��9T��hl�6�g��U�J���Gi�O	Y�Sc��?��J���͋+��,�jy=	@*<�_&��^)Q���s�����n�
 
���2�ej��5��|����:��?KN5��XZՀ�Ö�&#����HRƾ]�aqn�Ta
MR��� e�;!��T.�p;q(��T�a��	�î4I����j6��_�	�0�Ii����89���_�[�	l4B�2�vt]n�ɑn��H�&ly��ʼX�ߏ����X��I�I�?j� ��v��P@����q�XlxVHYEB    1d01     a207����0�O�H��u�W<�B���R!h��ôoĨ�U
'K��瘒b4��׶]x}��E��iM��;9+��)�Z����Ԭe�05�i͋���H&�0�1��8@�o��9c"#�@��J�>�g-CҘ��̄�����Q��FO�2�ub���y�4K���V�#�@��|��<�C����Z�<n��P0��%�_�P<G�͟��l�#�ќan#�Bh�n��!�W}�g�W��5�<jT�����D���a5�Ǜ��FU��G����b����<إp����f�b]F��R�~Ueʫ�S�M��^�O�ˁ�)0
�0�=�W�"��Ԭ8h�Oۆ\������#��$=� ��ރVI�]G��|�3� )�Wt��}��c���c��/6"i�<��[�[0��w�֙�J�B������e����7n�|?���nK��N�۲~�gE0@hPS$C;�4�án���v� �h\�`$�i�7
>���D��Σ�M��~��W����
c�o�:(/�9C���T��{�[O�lY�lȢJXRn���e����GĈ����9���/Wk*|���V�?E��?�i۶�}���B��y:]�~�4M�1oGs�����s)��0>��A����������� K��DH1����H\��U �W��.���6U̮��O�i���(�6)�(��[}R��c�Pw�Dp�ġc�C��=lG�Μ:�h��Wmv���44�.܀�S����,�=��f���{Q?`����_���`7H�nji��
(���ر�w*�U�y�P���QI�9����~D�����HH֕	�U�R�GP(�|9�@Q��x���������F�<�*�E��=y��˼�Ǯ�Ǚ��c��ĵ����
��'(��  �p���F�BM�ㅧ3\��n�:	����4Jx��J��z��xi{��/ظ�)�e�@���B9�ї�~��<)C��Z0��Bo����q��.�+����DTE��]�ϔJ��6`m��&-�*�aw&|mBB�/�A��?Za*Fػ���I�8�������5v���vgp�1�'�XT�N8]RT~݊�Cד��Ve�?�r�j�Cʤ"eǪ]��۰���LF��]l��	����(	���<�A�&���Y����*�ؑ9$F��܇^_�7.	�T�z�M� ��I_�845,�ˍ��PY��X8����g�ďe�@��B�!�{xdJ�s�*�+.����f$��~��p�"�v�?S<A�t=�=��\�9����5���ѵ�� ����l�3�{$��蝹���vFٽ�)آ�7��W������c�n}4Y���Q|>}t�z�zq^�m�H�
��Ld�M���ڊ��p`a�O��l �'-�����d.o��D�+�y&a~�\�/���ZV���"P�I�^Ƴ�E��7S�W1�i)#��#V'=P�g���h��<$N-c�a��e+�5�(a�M"���?�����Es&�2e�6'�{�����f��|�яV��!�K��Y��aN�O��P�h�a*/êO�����a���`SX76�W�k��ٲ�?'Hc�G#�>1v�T�thAM
��AgG%YӢ[���J�$���DV� �,�� ���;�}�2���P�T@F��z����/+V~z��f��h�Up���%��`M�C�.��h'�o �5���)k�y>21�+�݄2�ﾫ9R�_��3�Wi[�@�V�u#n���J��%�Ͳ�I�^Vh<����(�3]��/b���y�<�JI.k P�Q��#�M�įc�f^$SY�)�)�S��R;�R��dɻ�������;`�K����]ٔo��"�]x�Y�ퟛI��[ۋ��2��'���;e�"g��t8��[�up�c|sp�*mW2�"s�G/+�,+�#EŔp<��‱�r!�D���.��i�s�e}_�G&$�cR�u���H��Č��,�h�$�|���%��� ^k�b�aXA���xN�Ã��˫sj1�U�V���l�]{���1��%�I����x����i���-���Lm^�%W0�u%�:�WW���B�2��^���7G}�R�c�Q��K���C����4��֒��{n�a��0~�̉�7��N�bD���� -��k��f��xdl]�U<E���IS�� 8.�E�ߧ���JL�@�,��_�Fz��	)sL�h�y��^�֌��J9�A��<=��hZo��f�t�V�!q��\I����u� ���k��kp�rC޽�9��.8;aI���XW$)����ϲ��N��Hr]�LMmO6�\��^�!	\�f�FD)bV�C�+�~�w"巇��R�k���ۂ6�̽�j�qFt��A=道���ϑ:�C����4�9��h�?�p)��2�*�z�fW��H���s�ʫ|��H^��3��`����v0� �"�	�H2�MZ��q�R�u����6E��Sp�韬h������o�<�|R