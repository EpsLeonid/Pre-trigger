XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����zXhOD�{�%�&�).�����wD.Y�Hфz�@bgUX�����k��Y$�m�}BC}�/u�����.�������*��r-~ul�?�	������g�)�:���?���x8�)^�_dC�h�o�v�>�%�V�O�����2���k;0]�\ç@��E���j�В!nP^��NV�\}�9PQ�[�'�2�Q&C�`_��4׃���wu�r����Ｓ��zPD^n
6�en3h���~�do�*�}�E�!7� Hs�`��� ̿��Ҿ]���_Lt�/�5���˓b.W�=�����t�OgR|gu�$p�����[�Ip��@3#f���*~��T���3~���h�j�����hՀI��ң)��ކ-H_�N�aXs�}
:�;��r��g�L���k9w��b	�ˎ�no|�K�C����gn�^�z�i�����ė�\&Dp�u)�X�j�ɞw�=�s�B^WQ%�w�9��1ݰ]-�e%rW��p�%a?P�5�Ҩ\V���"�^R��  �7�C'�NCJ;A�ۮ�8�ث��/c���e�_l�Is�R_&�l�}�2vU���[U쎎�_`�.(Xe����5�!��e��B���_���0t��=c�G�za�E�@8�����%�iK�􀗸2�}m��\1<3ZW�g8h@���B6`TI���G��42~�hO~r$�!l>6U����a��.6"c�ƥ��íC��s��U(������XlxVHYEB    2327     a90�n���RPH^^�?�ഊ��rђ�q�!�, ���Ϻ�}
��0YG�t����''F��.Ww����;���_�(M��L�u��&e;��zGQ����CpY�5%���iPQ���ϟ"����f�Zl��6�f�6N_X�en�����l_��S�W0��7�*J�ݰ�^dX;DQ�
['�c��OM[��1̸aH1-�����>F7% P%�DX�}�}z�p�
�T��ǵ��.�S�[Ih�_�3����0� �p���d(myYZ(S��DR�G\�k��O��ȝ=p�p.ݐ��{�~k��0�k�g�^8O�ߜ�2�H����6+�}̩t�(1K�	!���E�g�x,�B@ǭ��`����G���s�#�h0�$���^�^"z)�6|���d}�"��C�Y��J��.���ў�C��� rSc��-�O�y��3Y#����G@7ė����Kf�����;\��7��G��R@�	���?�� ���B ʎp/��Xڬ1U�����<��r������䠠[��ѹ�M���eTzs��朇s�P:[%���I-�jI����F��4I�5RƸ�Ʈ����5��(@X
���p:�dQ�3�s��� !N?EmNރ��aa�[����y�^��-�yk��'L�rjڪ��#���5�E��<�=���%KR.��e���,oH����+��N#@l�/ˎK�]�s�An���Z��n�L����P�o�e5D��䱊�0�a�P� g�~��̪�	�����\!���������U^��D5�R�X��D�����q��� �n�Cr��K�437|/܀,�����x�'��W�Py��R���@��/�<����-�;q���M���6jJJR#2��\��ᎆ��6"��9:N�������@n+^�����h���Z�D��M���un
�;�1��r4߾Ѳ�'�x [:�M&,�������\Zap�-�q̸��,����'uw��؞��Y���a�M�D��F��sÞ��V�&tZ�è�[nJl���~�B��hZ ��c����ܪF��q�1)�B�'T����t(��Tҟ��\�"�-X�>6l}wh��IG.�W����س�/MK�;1����*�!�>�*��hÁ���r��z�����}<��H���"9.U������ձ�0`BM�@��Ȇ�FOC��V�G��:����/��"#�`}H�<��.xoz�J	)0�/��$4)�\�!�5�����H�1��q��8ME�Gch	NR�1]ݹ��J��u����w]���'b�]��oF������!W��BC��/�[a��HtT�PjΡud�R^����~������tq�Np._|��s,�G3�e�y�u�cʼ,^�RdS4_�&�Pk�My�����2P2޿��~sr�E�F���6���oQ���X�
P�`-�L�2;���+&�X~�=+N�hX�x�5��2�0@Q��q��_+�p+���8�����_#��w;2�`I���o,W*��N����$,1|I��5�{3��M]6:a)�������;Mp�;!�@��bPof򬠄�u�S��l�{�@dEH@�6�K��Bp�A������{����TH�⤨;l(H(�-Lh���&����r]ڈq7-��>� ��Y��EY�Q��J4ǂ�p\뚀*}��9�{bV����G�i�z�Cse	7��兜����L&�����r����1֊%N��H��ү��Z�G��N|ZsF�$Xy*q��ۄ�T�VC&r��6mRL�����8
�j65��ȸ���>���ʯq�}K���O�LM�C	ϸэ<��Ǣg��Q�z��ꊤ�F���?̓���_�;مW����R� ���󮭷���Vu� [�_����I��U�	�o ���费���>���]�ɼ��+������kgI���iDu�s󸰀ߘg�MТ���5��0p!��ęvNm��S���3�X0<�@�&�˷UK7]QÃ���<��d�3F؛�������a'�L�/B"A��KYzi���Z���(��K`���O��1 ۄ_&��-�*�=-{���9��@m6�6�.e��_趠���1��5�h�6�����f�Po���,_�D������ƃ#�nĊ ���h����20�ƛx:om���.pN4P�L�A�d	�LU>:Xp>���'M�{Ү��pK��(쌚������<U�4�ϓžY���Q�n�<���9��!ܱ:�����'�@�l���.�u��M�^�P�4��LM���Kv/�,|)��/���ϢCDk��N�%y-�8jh��p��'�x��x��d��(�-(
��#zZ�<�q����(^���\��,
�iM��d��G=w�`O��r���I�+��*��zTӕ�Z.[X�Q�/r�X(p���s�T��E$�� ���.�וE�0���No�'X�����U��\ED5�ZJ]
}	8Fj}ܔ��Y� ��@�֮&C@���Ω [��m|2�D�T���T��ۢ����EC+��/d u\և�7��w�d�2�͞��q��4���1��S�j��s�ij @i)��R�h9a��ݱ��