XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���d���]!_��Z+O=�	��)6��#5��V3{INl]�W�gE��%����ɣ�W��u8<��K��4G<��\��8�%�i��N���t��Y���5�a���|�l�ɏ��u�Hƌ����P.�|��c����C�tkq�H_f����%��P���u���tM@z�x�ߜ�`G�Za�//����q����d��Z �8��V� (�#����P�
�]_@ѝ,�lsYwҹ)�<j�O\*�w{;�QN�Y���@���x��r�EF��҆��@1*���TT-�\�n�J<�a�!�dnnX(~m�@ȑ/@f,Aۼs�Q�Z̼R��G����-���(m�ӓS�M���.?�v4�����[�`Q����GȰ탕^w�C�*IR&^���$�Z�{����D��T�c�θ���Im6�z|-2�L7��X#9 ߛ>��*q��*v���j��ֶʡh�]��6�&Υ�$��!+����Ilz3�2-��@�޳���!t�Yv������1J��V01�{9S
ZZG��G��C�� Y�ä��
�`jt5\j��j� �B{TTG�����Ʋ���m��OU;�ϸBoD�զH��gCd�xq5��)�\�Ɠ��a�A2|��:R��\�q�]����^y��B�'#o����^'�N��3dY�tc��۳ķ���������3˛g��c`�݉��.�9Լ�}9��Q%���3j�BzE� ��T�5e_�*�Y�XlxVHYEB    159e     7e0I#%:B0綣>hy�p�ɧ��"n�tB���~؋(��K�"M�<7؊i��|��N��h�J�L�A�]/�Y��s�������t`ɝ��	�r��x���
����W����$3�E<K�Q��I�*>`��%��{�+���Y�}zr8�p��e�!ϫe��9��p_�	5�O:��v��q��p�T�j�Zz6喇o2��@$U�i�Q�}8���L$c�֘z�h^ �G�mN��!-ǇXw7��pFdF7�-*g�{
γ������h�X��7n��c'M�����I���"�}���c�a��`���M@�D��Tq`�Ҽ�\�I+�C���R I{h�#�����L!"z�eG\b��P��l]T�v@�ˢ��Rt�|6�\�\W�tJ'@�BP�Ւ�3:3ł$S�vS=��c��&�}���ED��u�Y�1.}@��'RԈ�y�l
��|�K��e�[ֶƼ���=R�JN��#���|3X���k������&>1b�<2�q�y��l�o/zF��HS3a�]��y��6��� ����ծfW����(\�y���m�b�R��`�@ٽ�n�ET��ڞ*�0�<F���l����i�c����[��N�W��՘�8�E��+r�� �d�I�F�_�;d�ʡ��g�|���C��:�mJp�ȴ׈�6~�j�cO�)��<�;�cSXv*�k��̏��-�>�Y위SA���C�(��!@�I�iy>7���zPu,��.Ġī/!Q�m���a9K��f�E��zX�:��4�v(��KP�����{?��� >i���ƭ����G|o�k�b�`���N�[�ޮ����4�|groOqxvwΆ��U|�!�8���:���ɽ���y�c̏��'�=|�Qt~�<�5�4�q�ͷ�@K�>
�f�UXI
ҭ@��f�{w`Sܼn�W\B�Є��G��F�m����F�	�,��k��%yl��N��i}��1(E�ńj�R̀ۉ3��+����h��3�B{�g�@�=�i�:v`_,�L(lqw���Rv�ps��7�}��B��y�4~��}X�^n����I��A��3@W�#��M'*+;gd�,���5�<��&DC+���������~�>/�P��=�t<2�6��)r�L-�P(�O-y�䚯%�l��ͪ��ώ4���FH����S_��A�c���fa��ފ�D=	#��v��^ r!�Y)c�{.e�lz�tQzy��#|Y7ߛ!��JЂ-i�jk�0h����_;H��2a�4/���K�D�ީ�L/�����C����g^[QSM��1�)WM�V|2���̕������MM�,vIN|"�1��)jbQs�:O !�/�ܖ�s�F�sF��`'��z�፲�pS~#�W�i�6a��9Ϧ�` p��G|]=Br�<�;#���M33��ސ��K_��|�!�6�t8~�|۹W*��JO�d��Q�-�-�`/�Xa�̏a�Y�C��%Y<~3.���04t�T}����Ml��,��$3�M�TxC>;L���̆�t�\'`�H�����4Ê�FP��,���ܩtl�%���
�*�O�t}�X�D�ޙ�΁ �N�^�����N���������k��ǒޥ��P��|�h?�{纳�`J�EM��Q&|sթ����A��~�qp��i|�'�d��$��WB�gl)= �*�Ԕe��L3�s�A��>��C�%�w�2�֐�����n&�%k����a�T��)��!ڟ�}c��� 2�`<�&A�z��=��B(5�jb���I�_��f}�,FFOm�mbm����]2`q�0�����,����Pu6ĸo񰶹G�:��\�e�n]7���X��(�L��ޔcp�uI�A�����`�t4����eE:zA�-�2��R=� ��wŤ�a����^nC���e@{_�D\�D���\��$f�+���&/