XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���p��;=_�zP����V�Z��>��]�l�W(!Z��P+j��D�b�_fK��^EA!U�,�oZ+�p	�#�}��O���K-�
c,K��a�ٕ"q#>��8�b&��{�)��H���Ρ|v^`�K��Ʌ��-�!�+ͦ��kͭ3�����F�G�=�֎��`s��ª*�kHN���/ρ 0����r�>|r�f-;L�O��nw�x^�KEvS����i��!$I�R�Ԩ�7�k%�ӡogt��k�K��h�Qo'�����}v����,��2�0;��v��X����eũ�+Yd9���&vf����=�53Grƛ�<��9Lt����|��D�����c�=�Gc��E������ߓ*�рT�=�������V�'��nUo͜�v	:E��X�5h�i�Zئ��Ov��]U2��.�ܾ�E�WY�/G
�������N�\�)��]�fˢ�3V�d,���m/��E���``U��B�po)9znB���;C��`"�9od��ڛXe�q�]l���k
Ϧ0;���$��@,�c	�^ �f�]���V��LBIl����[��<��b-T[R<�c�B(o��TR8�<���*R-�ue��8��K�1��_�z���weD+�v�45��[§V�g-��.�(v�j��qA\!rLHB2P|�(��q�/!������k%��v����m��1�yNm�y>���I����7q���jsv��[3����*�Z�t-�)��5����=e�� XlxVHYEB    1661     760O�>D,{�/�?k��>;~��5`d�i�!�/���*DKF�6�����u��y���SM��jܥKfa.��V;�}�\������J� ��3�YGV>F9���)䣮#�;����^�U3����PB	Hu���S�6i�5b��ڇ���(��)��l>,�v�üV2�ϗ�B����ŭ��c�v2�J��t(  ���,��m���c�h&�=5�Dcxg��8��F,�T�q�2?�=Ⱥ
Qy�0m����<D�;��#���R��$�!�p��dr���e�ZU�mP9��4����I��&���M�˃����	�|g��[��P���ܴ��}�Vk.b
a�{M��~����x�ro����` j؟K�,�D��v.I#�4��r�p��J�z��?�2�.ڒo@��Ԫ/9��T�X�}�����D)�>�_,����}|��#Bkp�_5l�=�je9�n���C�g��1+�
���� }v� 47��ʼ�Hs��y#]ϫ��db�ߌ��jUock�ei�oa�3�k/o��a0���P�nHu��5�X�l7�7�ܹo�0N|�#U�h4���Z�����]Fn�WOO&�[0��0�h��(�w�8m���ݜ�)5�����r���ݴ�bنak����r>��Txڝ%�iY�n�*�b햛̙��Av�b��۠?��:��Az@K(�;)C�d���\
�ڢC��}A�%Q�q��E������+�4�Wh^���+��ƖꤥC��0�������`s�_B�~��uH���@�b��-��$^���� �8-��5����ڝ�$��?]!����k��'��z���;;aX�lO	�Pv�����ǳ�f�d�+R�ͩ�i0S��l԰K��v�
.ׁ�ToSJO���D�7��7�ѹʃ"W7.>s�8���9����S:�8�gA#����c�aM�B'��R�Y m"�d>���qQ����	Ȯr��^UF���n�6�V�����24��b��F��NK��X��5j�p�-�Г�Ix4]2*�wl���+��s�[�c�i��wFB�R�| �<b�8Y2��ДV���� ���qAqqQP�ǖ���8׫m��A>���ֺkByr�c7�^�������6������{�#,������,�ٮ�n +v�rc�Z���+_:�9�E_+�5��p ���i�S�U���U�|.�.
-�%�O��R£u�[�[_i72������(r�(Ť�,��h֝�������
%�_6�ꀭ�W��@7~�P����kY��~$!��D{��1�������7�_ӗ����*6�9	�ɖƭ�}椲w�a��=�
6=uȴ(�Gd�i^F���*KN�v0��� ���Ě�T0!���E/��ɐ�-�����B�`�Ҙ��I����GA�ʹ8*�B�����w�Xf��7���������A��;B"�Qu�	�T��
)��Mɐor@�������zZ|A*�:�D���;�W3�Eb�T��!Ev4PR��E񝻪@k��9����u�s~���
 ���s���2��U-��%ҷ���[6TkD&�&�߂��|�A�û����ż}�x��砭�m<��������
UW�`7�"�PͶ>a=(����Tֹ��PԞ>B�Sξ,D9p�0r:��� "(��@��t����h��ot^t}3�����d{��OȅWes;�xs*��͂��|��x��:,����>��oBf��]5Q��a1�ؐ3����m�����
l�BWy���Ԇ�v�d�}3�^;�^�p��gP�R�9���;�t�!�3]�g,�?�=��pr��u;