XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���m8~PN`�v���o	7��
��q 0�j��a�ܚ��<�^-�{3d�"�?�Ȥ�#U��b�
�:�ك(�����.��v�>�wk�tm�4�Wm0F�>�2ox�®*롶"H���KsI�W!qq���4�����ɣ��������_t?dfo{�����cJ?�A���oW�p��Q'���k��s�p�����f���L2M��5wL�`曪�Up����1Kk&)ǰ�Q���4�˷����l�O�
ׯ�~e��L���Z$����dc�p7ڤ����NWF~�\���}�֌����qF&��-�C��BG�r�^[�����:Nc�{9�Z��W�J�������{T�������q���^F\[�5��pĪE�&EEr�k�t�� �0zSǈ�Um ���.��SG�M�6i�?����H��"�f>���b~�m�����|;Ģ쳤)�*�24|>����+���>#�p]�`���Ƞ�6J�x���|a5�����G;��:7��4��n�<À�`߭D~�#��oO�)��Y�r�!����b��A�����X�X����e��{��?[���3�f��X�e#=�g}����ݼe	�0�Y�d��>\�	տ\3��l��]��W�;�K��п��f��|y�j��X�l�����ls����`���(Jg�d]A*�8B�x-�a�sя�+m�C��a�B6��͙[�Կ3N�nH�p	^�ʒjP��y����*��sE�&�XlxVHYEB    5fd1    17101�! �����]�*�d*T�c��f�W�����;�j��{5F��J�]���~z�x���D#<����V��o�2lb�I�a�_�Z���J�J�G5���U���W@�C�-2x��VY�7�{pL���ԉ*V���.���x*�E�!j��r��b�tɯ[:�o�r��vi��%�B�d^`٪�K����@;+����<�Τrg8����k���������ք@�Ù�2�fj���Y�������!��f���Y�W��B�k�	�b�8������
��� e�S�)��F���T�������V�1zi�S��_&
Q`�BQr��+�כlg��&(ͼ꣱x�P���h^��u���Զ3���Z��8�
�yc�}��B��dx�C;�f:i�����<�(h�|�8h�Ƀ�TIC��D�|�֑�{�F�*�ċv�^��d[���.��}�n��qr��uX��o�c�r��2*ڋ��_�9��Ǭ�89��wgJ�)��7�ן9�e�`x�
���ިǌ�+e��X cr�D���U�fq�Lf�0��,�Q%!_mf�0��*&�˿�����!ܸ>&���T��=�5�HۼaNw�\MzS��3aBA�=���ܿ�!/{t������_��������}�����O)"N6[DX�sS�V�	d�½����^���FV�Y,�R���<t��6��Z�՘���~M袣��w����JזԬ�d6�sK�9Z: ���2OU`�ݯ���'ֹ�y����U;��˩���rD��#H0��Bf��|2'�-�b[>F e�q���|�N���zL��vz��{���s
�)/���,�ݱ����lW�U�+@�� ��.	{Nb�fy��@|͟�^v��|P��y<�i|%{)��Upu٨����>�ף+�K�p	��Z2m` ��=��b�.n3ߵc{�f��v�l��M�(�{�h^a��W�8W����%{x]��≠,?(���p�p ��uƱuDW]��gYu�o/4�+�2d�Vi̥(ʡ.a0hY��m��9�Gۚ���b��j�Dޱ.��֙<D����gQ�#
���#� ����W2���=^m����9bGûO2ƾc�&� �o	b�>��D���
o����,Y�b��'������Y�ԱT[B8o�c�Þ�Q��x�w�L���������l4����cدz�<�����ҵl�p�8�ob= ��|�g����ɓ=��J�����S��y����*��.���I��Ԑ-�s16�NS<FǪ)p���w>f+5X��%(6ҋ5n�=�A�$�w1cU� C���q���d���RSp�inc!��׻�d�;���Y�V�uB�2��]��C^�ā�;3u��6!�H����\�uG���jR>`���/���L��^p�|"�#�k�/B����_e����9�͎�"�~��4<��iq	�'�Y���x��r�H2���`���ch�[<�<�lOU0x#��������}�8�8�}�<����F�?+T��"����P�)��xn�+�!�q����/R�0r`�;*�%m�>JRW���W���H��Ti�T$��t�k��ug�zeXz·���͌��N�o<y�N�i1�Jk
-�]4	��G�C�G�t�V���z�b
���+��3�#BG9�H|�`˴��{V:!��NLL�[/�\ U��ޟ)�?��b�DR$����XB&\7�����]�QQ��F�֩�ԭ��hհ���^Z�u�騬�;Ժ!�V��2\����o��˳�C���)�t�9?0�~7�D:ž��l>vM�W�GU�e�[<�W�Sm�÷_����������Oq���$$<]�-м⊶�^^+���z�����l�>�<���W�_â��rM�4��å$���T���z���MZ�w':�$Gw�6� ��b����6ű�����3��G_ܘ=[�rz��[���J�rw4��Q4��nT�aFQ��F�)bb�J���ц.1��f��0[P�0�Z�Dt��w��0��M��:�PW�i��~H��DR��Z��wd.����h�q�ࡓ_C��� v ���6h���j�|p/��i���XE���iP���ns�ʪ{k�6��sɗ&����Ea+X�a��(��AQ�y���!?.��5�;���Vb���b+�g�]4��8�?/����9c�ܛ� Vfz-N=�l��U$��SkRNkȻK���N�nwb	S��tc)��!vW�-m�F�P��=�����	��s����P ��=2j����v�I�KT���_�(�_��oԼ���r�w��FMQ"�:���ȧ۱y'SѦ)��:W9�P��r���/'T�ӓ�Y����R�p�sF��J�7I��!�^�ӀC���G�\�$����.2g��Ja�EO6Uu |E{+ͧ��+Ё*dS����P�"�Sm�"Z�`��k�) �����IQ I�~�9Gz<�\�C��x���R���L���S(�&Q����|+��2Đ�K�ן5�ԬLk�������!z���[��D0��x�y���qi����N�E��,I@\Կ�H���#���1�c���3�r}�T"�lg\2���� ��]��P��P-̣�?�4�*bl3TL�c7���'���`f��o4Զ���?7t��/��J��l5�>�b|��w��@\�ڥ�aٔ�orI`2�1�s�D��P�@oZ�V����3�)$�� "֓���������!3U�Tw�-�p�ǑbB�\��?��{�ɡ�i���˳�o�Y-'!M���b0'Bm��J�[<���^&��!�����W�_�l���{�ꛔ��>��{�
�P�dZ������T�������,y�ܮ�S�y�{��7)̗k"C��71�N����gD��nqf�� r&����	K��<�KlЧtW^��(M���l�-wئ���'��9����h>Ņv�����/y��{#q4�ǵ�@a�W!� �I��0�&I�E����TDNg�B���Bzv�5_�C��M`�  [Qza�mV�gw�1b��b^�o��Ԫ/l#zW?�B���TOL�!�V~Bí$-�bU�R�E����I;۷�W�����N�����U���X�Z��)T����_F�F�.XoN�#��T3=!@N����[�2PhB�԰:��4#��� ��ݷjX��`�%�j��B�З��l��
��koe��,�
@E��;�����B��� 5�S�>���C�}@A�D�P��6�-JCv�s�O�0؊�w�g���Ƥ�n!�:S-#~���b��4<�%�N�'��r���C��^DeC2fN�hqo��R��R 6��N;�	� :��o�w�;�0��ǐŦ�Y��e����Z���rK���Jn���`}�䫆I�c��A�r�X�1M�	Sܛ��z�Щuĉ�>��ǲ�A3�Y���y�q�N�q��89K�y���|6�Y��+�ucP�r���C��K���fa�W㜟i����'9�xc�z5t��WL��Q{���:�Z�	FvCX!�39:�Wb����J��$
�BU����_=jԐ��n����%�,���H ���-��d����b/�ЭIo�ă���e0J��j��O���gc�v���1djHk�>��P	�T3	,<�t�W�l�l�V~�l�-�TNBS�$%n!��ڦd���*P�&��.��k���Jqq5��u^�,�lV.���r�ND�#���(*|_�mI��4����ȴ?��,|@���]Bx�J��^�K�⊛��w�`���T�Иr���gk�2^��̎Y�K&hEE�\�:�\$u�e���5��e0.��XMHE�+�\�]�7B��c��/��F��OE!>�F�G)��Kp�N�c�U;g���ҿP'&���)�>!kRj����M^�uR�?ɗW�<}��v�Қ~�YA	���u;�3�y|bP�R�	�Wzp���%I�f�p�M���� RV�O���m�d��2�"�?�r�j<�d@���iX�^t���Uy�%+�̡�tᢹx��5X��h�E��{!�'O���)-�x�oB�Q�Ļ���'�q+�M�h�2�����9�r~�(����I�fM�B�k��|��p5��V=vc� N2�@4�@/L%�BA�w�|ow���ǜ˕[Ϧ�@	L^�������|C���*n�=�Kw2�4�_�Eކd�����OF;��.Zh՚� �?��9 ��o�`�8]T��ru�ݿ�0���C�>a����H�Z@y���B��'B�,��E���N���'�����5_�V����y�E�&⭬1�B���aFs2���A>n����TT��A �?�pHÜ����|�*_�QF; �::'��/6O��~�(��.p?6�E'P.�Wl�5rR�rHD�a�P�̎�qω����$	q��':�4jh�@�$Yܑ1���?l(y�l5M?�ȃ΃^�1b��2�`��:�޲04�ٯ���m������|����Y�{���U�t1�WR84���Ygր�]�֛��T>�@�x
�f~��A?�PM)�-4>�$�R�|3j~��&��w̽��������g~��SRd�YN�-����wm �N]:����~ޅ䕋�+�[�,�-֤o�?p*�v���ׂ�"�����X�!�M�7 ��۳�;8¨a\�O0�Iq�`]i�v������a�zA� �n]�!&ǘ��뢛	�@�t�	te��ʮU7@~G�Ǔ�f�>-~�4?��VSA�eC*�,��+�o����o,d/.n�LkٔeS D�Ws�cc����^�L �w"�!KZ������T�1��[�H%e!��R����
��"���W��w}��������/%����3��>Gqn*o[;�o*��,�~@+y��k�A�@�,ַ��*�<�â�Ύ�P_Y���W����5S���H���Ծ�k;N���]�A��b�z`U�~��Y�V��9�X��+-����cptӪ�g�Y���w��i�Q������]Uш����ux�qz3&eԅ��N�N28�Qe���BtE�N-�=���)c��P�֦8:1|R'N@c�>5D�oBs8����\r�|_���	
��&&X��y��eMI�+BCiK�J=�P�!Rگ!�TQ9w�)K
Yޡ%���r��FaC�~�"���aMvwuS.O��p+�8�Q�d��[� ��j�Qĕ�4���V"��7r�����=���r���׺X%L�"�EJ�5���u��y���"&>�hw_S�1u�솟#������4X��! ���T��]����``���G���އ����>+����GP�j9�"OHZ�4}��£Fg*	�8�Y����`*�蠢��!����dĠ`.x(�s�����T��ZY��Z���F[�[�:/�$L�r��1��9Wͥg���+=��)y��|�q�@�۩[<����6HI���ԡx[#�q��A���� p����%x�6�2l�5�N�,h[7�awKy�YZ��n�9�5��4����� ��)��n[���ς2�)�k�m^8�ڷ��i �49x��ڈ�sL2���Ѹ�!�����Q��4!�v&�
�S)�f�O:_���j��.����E�k�LJ{��	�}@�b�����@z�W�`���cf��a�^}I��s1Mr��v�̋8@��#��F4!���c�c��T�'�2���v