XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����ŗG ���8��K���d-�F|of��|-k�'1E���{��@��-�\��C�#��� ��{tAW�G#����V�V��~-�K�;X��Y�;�����VmgW4��4�6L�@FM���o��//�)���!v�S��$	��kj&���j�5�G=��M�0���`��05�ӗ��E���7��o�Sh�R�!"��b���䱿{�a�����=d���H(�$��de�8m�]��u�J�N����#'�)�ss��x���L�R�s�� v��$R��.�"NM��@�(�6�Y��_(?J���J��S��Vj�C�����1�z���ݕ�J�) 7�c#��K�����l~j`��J��-�A�Z������|m��?���)�I�O��ܚ]��k�F�1	/��TX E�g�iu��Q��ȼ�}�;u���_eN3�祠�KD͝�9��K䷍�M��L\�Ë[#%N�;e>{��躋J�~�i�� ����$�"��*ה�^�S>�*d�J]��l����ܴ>K�N�w����k�Sj�Ϩ��Lz袖����R�*���rѓd6�(��N´�SmO�:�V[vo��X�|5��2Y�כ� �eNj�@qM��d���=܆p�K�[�DL]�oiDm��T��K��K�RP���)/@U^*�+�[�)�3Mc��
���7�W\�N�r��x\�����:���"(�ʡ��uO���g��b�7O�ϓ��mˤ˴Xv2��{
^�~iXlxVHYEB    5658    14e0V��5֔�݈dA��&�;7�#=��Wĕl
ľ{*��}J�Y+9�e-�p�� �ܟ"����;� �u�	������ÎG��8��Ӿ�'h � ����G�?��&KH�a��������^]=ܧ��8�n����^� ,/������� �����!9��|N�%�@���5������!�Rpha��r��Oh�
�U�%�0���7��M��M�,*��dU5���F�ܛOF�zlNl8ik�\_��ǧ`{���y��d�vQ],@�=Š�8��B!D��k2�f�+�0`�j�~�����>	��cܪ�W6J��p���t)z��w�n��|�?f-�C�
�74 ԓ'2S>H m���&y�:a�q��g��V�!sm�T�s�ҋ��kأ�!�Ӯ�����/��EVfy�!�6ʗRP�'s�;C$$A_y/�Bk$U���E����3�����n�`���ѹbd�HYg����?#�k^MR��"���3/
��d���M��̲V��1^g���PܩT��>��j��WO�}�(B�W�j$K��3yu�D�U�a�a]7$L�ݸ��q���r'�O£�E�RZ�	�_m�}q^�6�>%����{),d$�zȴ���	�M��X�ɷ�[���|2��lҢ��r*�oX�����Cs3��iC<�=�@eS|Ū���j��W�����۠\jS`R��3i�"��L�޺%���K�����u�q�\����h��-�06s[-By_!F���r�EcA^H��W�h��u���w�sX"D���`�����X3�<`��]@�+,�mOc^Q�օc��Q����k��_u���:��%b��;#�IrM�2m+J�s*��2��˾/H�!Z	FNz���p�}�`F����,��@kk#4ȿ��W��h�>��� y�d\;���,
��&(��*�[��X��b|�!��E� ��_/�@����A5:m�	l���Ś$=���E�o_-�v�zf���	��a��v��y��~��%p�UI��"в����Ӕ�����n#-�!��C�J�/�Q_�\�H?�$O��T4��y�\jP�4J�L�mt'ɮ|݂W;"�gF�@v�ϐܳw'��l<��{;z�.q�b�t8�@>��j8�4�C���R2
�-T���  �8\$0��*浢�Rki}����w��3_����*�)`��7���ľ�@�n.5aV�@�E�E���s�=����@����4uВ)�3�X�J�
)�c���;���{��Q�Q4ZH��**�C�2�[���p�`8���)�7M� )���lt��
��O��ƣ� �h�d}��M9]�UL�9�+`a��yb�����<U
j��·h_@�2�x��ԢsR�ybUy��7d�Ā�FD���1�2�V�٣�em�:�U�����l�>$��,H*�@T3��9���j�!u���j�C�9�s�\����_"Kb�m�U
���!omGСS�_�
��Q M�����w��I�Zi&�GS��6	+�ӷ�{�w�'��uWbB���1YCB�jҰ?�/Ξ4�zΛ�\��>�.i���,èB�?W�o5�����h`��Lu�~�'3`fq��FLA���cq���~W��6��#/�����0WKu������s��`�"�y�d�o23����c��T;ŗ�ʯ�~c���;V������oI��N��q�Q
��FO��@� �OV��,6�aq�Hb�8I��M�cG����c���!��d��_���B�q��'}IPo<�^0n��Q�vK�߰M����L�r�)��i��I�\ ��|��U�Q�4�+O���T4��[[y�Ӥae��DDs��s��`�v( N3�]��'E�������*�Ե��=���~u�_I��A	r��"��N�
xg$�;I9�C�����Uej��[^6Q)�IH���{�3��W節I�H��=�pdI4t"P��j~{�������I�򏺲�%u�O/]Fp;����Д������ߐ��6k�t��w�}v��z�"۞�Y7�X�%i�L�{
����E��/�G��O��,�|�K�D;kZ4�	�� (03��.o&��.����w`���X��Jv;r�`漐�u1�C��C��,M�u՘�	�Y2>�oo�Hl1�� R�j��]r[��4��P���]�Yw���9�.ȹ��.0R���YV�������:���r9�I�
!��W�}��gt�-#��VϖC�B���y�&�����/B���z�<B�	o夰�[�z�)v4�#�ƛ�?)5�b2��a�-�%��v�.2��o�o��s�i�?�S7�U�ڹ�(3�k�R�0�K����q��24��<E�����>�|7�Ԅ�㍱֦#������Q�Rv�¼.f!>�N�h+s��GM\�l/Y_q����Z�h���j~	u<5��)��(]A�lq�C���d�5�����P�	�g+=08�I~C��i�<�����А./#���,�*�s�n������-Or�^�g��|�d���\M�k[D8�~"���?�_%�d��|�,�ƾO�}2�R4[��V:�_�s"*p ��"v��OU���*��B���c���Ϡ�rY*G����A{����(�,}E�ߖ#�'��� �g��3˕���0jFU/|$�����7���U�o)�;sm@��i�J&Ud�Қ�z|��z"�N��Ng"��EaG�
�`̆�b$X7��$��2Nu�U���ZW5��d*��>��5��r�Y��AY��p�E:q��{	���?6�v�3�J(�BF���Uw�~I�f��n�MKՏ_C��ClN��y�%��!�t�Ǻ@�d@�D;I�I��}gZ=y���!�f��s@1+�3���}t��y��@a�?{��4�N�c���h�Q�x�^�������	|>D�3��G���ǵ������PۧW�A��� oW�}ME�tJ�H�[b��]+oU����S�v�FoT�x
��OK�T��݋�7�n�h�s���p 	&2U�d��� Z"
�(_7k��M�� ���� @�hn����Nd�����[�}%�IO �ߙ�◴<
�
����� $�@�i�Y�Q��Z����۟�7V�U:��q�󂦨�Ń�Z��>6��5:�u����u�pOw;͉B��S�[��HY
��wf��@u��SY���Y��g�M(�7�E|�������v@y6%���iX�޿��� ���	-�(�-'�h�fv�nJ���7}��$DbH��lx$�D� �M��G_��ve[Q�4{� ��>� �������7�����_����h$����U�3h$ZEǱ����WnvQ��.t&(���n�C�_�^P����ke�����#�"��˞�t�9qs��x�?9AB�/�k��Sn.���Q Ϙ]�V�(K�QD�m� ��j��m�`䉏�f�EIi��p�K�r����R�Q�&\�S*p,�f�¤W�>n&�w�(��x?Z��/��"Y��uX)�]&�͆������:)�_�� ����%<�[dF�?DTsg?��۴B��%r3҃~�J�����kʳ?�T��>b�a���S���t������$��u�L��g��ƽ��6�ar��b,��*���ߢ�Y!��j���;
_�PGö*W�j�1[$�����겨��B�/`b^~��̭�޴�O�]���<������	W8y�j�f(��A��z\�Mw$jy�w����Eh��]x������!�d؎l�qx��U1�s��d�DˌS�d���,�iT��t�^-�^.�(?Ƞ�X�#��=���D�%�z���Iy��%7��G�~�u��Vٯ�>rx�E\�����R�ݮ�&ρI���c���ȑ���0�I�w��]@����i;K/�􏿤HK�����g|��-"߰�=˛��b'��c���?�|�b�tqH�^��`�X�7������ c���SC \��]<��j��L�f����Ϊw ���~�tA����Z
���H�;l�_���j�����u�Ds�X2J(T9�t�·z��A!�g����-Tʿ�g�y��B4���(�u�~ﻋ:�tj���ARZCH��TK��Y�r��H ЌJ��J:G�}��������a��f;��������挲����.v���wH��W:�!ec�0-n��i;u	�dq(�,���M��[پI���?8��9uX5�ǎj��1���F��-)BT�g5J ؠ��J#��מ6K����Ⱥ�O<���N�� �]"����+���f}GV|�[����MⳘ�1�I 2d�wF�$pid]_�)3z�"�P���n�`���6���d:Y�H�v�0��F�m���s(����}����q�uV�gj���>$��4�S2"׭�;�~��{��i��f�������i�xS����\����9>��>s�Ӓ�����y���7�S�'?s�!5��q���p�3M�A�Z�6Om��	�j[;E��C��d��u�:�Ҵ
;�$��,�I%���\�+���������T��͂!���o��/�����7�aE��G�n��}ɾ�X��2��������R8����o+ǁPA�6����3`�40SeYz�"͕#G�]��<}I� =�\��0��Q�h��P��q@@�T���Zh�Ƒ��� >KS��A���X�;�\ds�{�I�s���;��@��(�h�˫QiU�����X������+��Xw�da�yr�+7�fqvpVרp]���Y~YAd&�%����֞p>���2b��d��c�\��n���;N(2ْ<X��?�������%�{*@�KB��1�cX�5jA�T��X�d�9��I98'��NXf�x��wU�&|�ޑ�>�	��઩�"iQY�v�)��is�~�^q�N��jB�43K�K�	̱�@^ďVJ����O���ί��u�:�bj�������4���R��{TO�o�Ӳ�stV��e���:�3#��7'��,�S*f�h9�>�(I��%u@�+�Gݤ?.��D������@�����c@�J�\�TWK�H)���]�W�'�M�:�������&%��86��/�Ur�N�-��Tڱք^Ҩ�54<�$C,�9�ޭAR��Bi�}i�9��� ��sq��.2�����aU|�D�V���Ӕ