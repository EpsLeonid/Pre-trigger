XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#הIC�[��v.eм\p/{��v�����k��ń�0l���:w'>�+Ī����8�]\b�JW���ձVH�h�h��%佂�_~�!��X��X͹�ꠍH�!P�!z59�,bR��-��O���7���V��'��w�'�k�c���¶�f�"�X6��u���&n�l�	���"fv���h����!�R���-!&Q�'��\X>��{[�o� �'.�p?�"D���>���ud���A��vw٬X�pdL}7�zP�����Q�gwT�G5���YȌC�Lǿ�`5@Jd���Y�r�
��|k^T���/��g�͟�[�.��6�4W4��N��#E!b��%!/��Bj�{MN*s�}�.4R�����/ya��U;�x[�	*w��l�T7�#m��%�����/{��� ��>a<�����BG�U�|���qDH(Q�>)�S�s�0E��a�r�֔�S�g�WX�/��E����Q��Y+�d��ui�LXfq�>mX
!1���di���C0��8A�-�}��oo�u*މI�,R���	���~���5�:~����^���:2R��B@�}�Wxx��P�L�,� �Ы�Y����H+D�'�0j[�|�n7i�Q�v>��.ϴe��NG}ѽ�2�1�:��>͒E�N�b�6�W��bT�Ka�u�޵u���G�Rh��:b���@�R��- �R�>X����
��>H�S��5?bi��n[����b���*XlxVHYEB    5571    1410h2����-����?�.R-+����|�|� ����3����O`��`��z|[N3BpMT�ӧL�7  9�u�;3*ӥ��\���3��G���7�����x�8�.�?�˟�1ŕ�Fv��#Y�� �[O.��ن�N6_�o`_
����1�i����������N��Y�d�1�M����1�rl�K89�ȧg��t�bz���u�G�N�$m`';E(��a@�f�NH4#@F��'��VF@�j�[�/����>d�2��/�������#�^~ؼ�=n
��^�߽@��<w}b^v_��}�����x��|���+l��;:�6K�\��oɻ�����40��L�:�F4��)���E0E���[�?ֹ����и	�,	WR���$���q���'$?h�-���u����1VV"���е+�(�x)�
�{}��t�G�持qO�?�`莀��8b���B���m��r�\<�ed�ɘx��z�ZϮH��Q�C�9����ŗ,�V��o�h�i��������������ar�ZP�O��_�ɝOoq�B{|Wk��R�Z��@s+�]�R,w'#��;(�W)f}4y=cw<5���5ͤC^���4�pk��vΨ�mA}_�ŗI��.�@!:��}!��(�sĝ۸/2v����W��.��u(��ۖ����|D��Q�Å-��}h�߾�²��9�Y��m��!H{�+�}���"��ڐ�r+瓖�
v�+J{��>H���� ��6�M*=tcG�����^�Ym��5��<��^�JL�����Ĩ�N����iǭ:�sq��� '��)�:�@&%]e[	P¬��
�#n�k�i�c Ox�8�{ܱ%����j�å�p~U08W���-n���b@4�60�*锚��`Y���i�{����M��.o��)���q��msK�����"X}���:,�m?Um)G�t4����+μ �@4Y���؋'��(l����5Ӣ���KJû�<g��˜�{��|��LB���'�B��M6ɑ�M��5���9�$�cyq�tΒ,�����-�A����~Ay<&�%���dW�WQ����3/�;gS��*�l�c���I T<�S�i(klL�
�ԯ�/s�	z��z^�V�X�ü8?�Ba� ���
�D_����Q�D�^�J����(a�2��*ĝ�����p:��}�:\��AO�OL�<�#�*4���}/�.eH.i[b��qr#$e)E\����:R����]�0���s�-��vT����.a�)���sv�J_�܍o_ש�h�^#*O��Z�x3�ԇ�r�K�E|2݀Œ�&z}T��Ax��k(�q�/�Տ��5���k�e�?�y&��e&�ZT-����^I�V�������5�D�����eR\�yw��~��Rv�&9�#��E{���������R���ui^�A�����+
�'c	wW!���Miq~8��z�5��|��vUBg߫���y\$~���5���XB ��`�B{���Z�HM!���q��Y
��K����b���I^��������ɆU&3��
/1m.�����#�e�A*�w���o�`�X3��v��PQ�t��2��Hb�˃0��9>���v�\�@��el62��c���|��GH��(v� {�Yj�+�
cVX��ȩ�u8���-��-�,�%�YN2q�-�)���l]6�:,��u�{��3�f��/����҆]�;�/M��a?�X�ږ�z�bjrc���ܻ|���!�N�dgl�9|��S������Un��f�j��ŖI�hހݕ��c0d`T���ȍ%����F.���T'iex����u�վ* �@�JWp<8�@�_�C�2&2ˎ�]!�:�o�֓%ϡY?Ad*�ý�5�����gn��U��N+}ַ(0�;.�	1�=׆�A-|kʂK[�{m�Sd��J���I��`����� �lTn��|��|5F��a�_�X�U�S�TFk^����Ld���Ad�>��a~��l�T�o��9�E�����b)����Q���~֋�W�Z9&Ј'��>����wC�V��}������¹7.j�i�N�DKY�R(�~�v���_�E|P�Sr�
�h��4g��:p�a:F�&2ux���+�%JR�=@�㛝�xJ�^���;�y ���ж��N��@<��kJ�Έ��}לӸ��е <�܀��K�����uP;���+7�ؐ]v5��b�A8���~���w�+���0�ۢӏF���������?��������m���xh���1�� ��{��u��~v�M�h�F�G������+rPX�8�m�֗u
����[V����C��W�pl�G���e���`6�����hW�d����o<������w�/<Ŗjƨg=�f���qpu�����۩b;��v�oz��_==�s���O�V��������`3W�]��
zWb?�i{�؊��J\.�*�Xn�E����;������ޞ[�Ռ�4A�X'�IKE�d$�2��,�ר�є(���,@ֶ?�ܒ$��+|F������߯���s;��.�5c�e��9�L�"��!�Ѩ+k\v0vNE�sF�x\0rΡ�l��3�j5V G����`Ԛ�e 	:��@�\'���"��oY=iЌ�DS;�Zw�V��D5���<��S#��t�~Lc`;�(y�&��/b����d�!�$��>�0��﷿�X����*վ����]U�8H�����H+�����9ziV�\]�c����i�A�/:0Bn*^��00�1��ЍZ����>�J�4�3�mF?h��w3��8�d�oC|�ʞ���ᤷ���,�*����������(=�˦�D�X���#�0)/Je6�FeHp����܅H�%�[��A<\�z.�0�;�E� ����tu�(�m��f�� q��ֺʨ�+�݃����+^�	���[�)b�pڽ�H pދ����̧U�����?[�N�x뿻�4_�Mޤ+��i��J��hv,�^��o~�0�SU�.L��D�DC�hph�ϵ�j?xc�R�!yI_7��H�����H�4�4�l�����(֥a
|�xi��-��
�O����U����RY���9�j�WPnN�T0�ڶ��OFNѡaO��[;l;�Ju�H#Q�a�h"��^�oq�����w4 ��x��D�&#n(�+Ɨ͞�-q���wvL������������v}?ފ������@����z��d����x$}�1Qm�4sA�̠e� ���G�σ;�����4�L�Q��z#@0�f���l
K7�4g<?�(�GH2��9�����0<���'��]�8�j���;D�~О3��#�\���O�_C�
jҮkBLW�yI�G�H�u�6�Q��
mr\w�q�x
����������tU�L���7�R@`�P� s�������7�1��г���x���yY�oݡԮ���Gdd�d�%�֩��3ЙO�M~��PF��`��S�ώ�����V�ȱ��r�N�8�s���1�8�Qϋ�ђ�ިk�}�5���e��y�t�1�4���Bn���<��,��,��p�1��لt�pA"�.Ӟ'�yTUC2�����oQ,e�*� ���0ɣ�? t��K��>\>�Q����ka�S�OC��kn�:(�ި#�y(�q�~��A�?�;�Ms�p��v?;�7$����8�3D��<�R-饫۰1�>z�.���D/Ѹ�Cx.	ͅuVp3h8?2��\T�nM��M�$�v/�.�0�����`E�8���˰�)�{�͈"���#�M�8��-��1gÖ ",qL�:��,.��K�Q�����̕�34A;B����Ϡ��%^B��
�-��V*�L�e��62��+ I�и�W����cxQZ/�=J�Ő|p<^e�e^�n�]�����
�;}͎�N7ᵳx��O(0��C�?썌�1���2I��g>���ӊ��F��L;��%l?�^��+���w`�5�r�Jy�-��3>�6*6g<p'e@CY�c�\^bD��	�J{�4-�Ȧ�����#��!�w����;CIY��f��] 	I����$Bw����RU>C@����?Ue=ц6,;ȫ���e>Q_�n|n���o��g~`���}e��5ғ���#�3�]�K}k�5��L�^��he���k[�����]��K�B`�'�@��Q^$�7j��WC׌�Ԧ^U�hj�	e8㜼9_[���^��iz�_z��"g�@���ɱ�+4\[�hL�i�!	�L��2�`�&t,z��*�!���R,T�u���T7.�e~����< @�nz*�>�����/V��M���LEQ���% ���1�oӭ6���:==���x63ڄ�� �Bq��R���\��W4XnڤH�rG�?�z0&�B����S���意�����l���"��J����^���,��¿����w�s�enC��<~�����!�w!U}-��&"@JUT莸�f�k���&��� �6x�4�8=BϪ�i."d%��	m�Pn%�F���WPHM������y�������t��>�8����VyVd�y�|�����vXE�Z�Y01����X�o{Q8Ǭ	}B�s�g�|�7�J�ZUI''G�Y��s�z��%��6��"��N��s�����/��E5ߗ:�):�׳���7�܄�$	Yw�k���c���5 C�UL�ͻ��o��=iq�%6�}Yh�d��	��3��G�N�,�_x���߈�����j�O��6<�Ѡ�.�w�4>�n����e��^��@�� �r��!9J�ч$V����ш����?2��k�G���y���0�g�L?ň����GyK����-6-y�]��?��b���&{��)_�2�)X�ھ>|2	w+#JXZl�`u�8�8�b�Y�u�Ovg8�4�7.6�ẏ1 �&��e�u�/���l|KmNDk�����v���\����@=