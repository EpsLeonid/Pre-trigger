XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Q��r� E�e;���m�[y"N�' �
����h�iBaC�~S%���IN��kI�F�(�@0��N�������摸�Z.���V�T���*}q5
��\A�[�j���� �s؜�=��,����8��d�kU��:7�@���,����������tK�2F��6{�w{s�
 ����`C�����l\�ڐ $�2� �d�_�!rmi��xw���`v�9��j�Z��4E��E�'�kHύLߝd�<Vn��L�����PCV�SӁ�����C��M�4�OtIfih���l��Â2��F��f�&�����(�O��h�λ�'�Olj�n]���%�V�<����E�0�Du�Z�50h��7|�]!;|Vq���p�xWs�F��8��O��n703�Ʊ���1�O���EK��3i6��k�\&Qv-<
�a˩`��30��̺��"���
?[[��`04�����cݨ-�1�<�7C�Q��ͱ�Z<�ZJU$˿�㴶ϋx�3�=�;���BfYk�4��GAjp����4{ p=1��-`@V�T�������_Mk��V����:C z�Y��[�������+��zEJ���{t�Pw�2P������MF�U���>��(�H*�a6`���î�ע��C���9=�Ϻ�D�\RGM?S��j;���b�EZ}G?a~۫,#��r���0°}N��Cŵ�B��1��E=�Y����if]����A�� ����_�*����5%XlxVHYEB    1d59     8c0XF���Ϻܞs3.{�/��d�f��F�#zgc{�_��0�S�A�J��9�'�xB!�-��RO�A�;��,���
ꧫd�:��}[̚/��]R2����
���;_�8�&�EO	/m���̽����E5I��|p0jGN�`� ��R��&̒��G�隓��u��@h, M�Bd�I׷�sMc7jX�^�!b�=$����j��	�NdՌB�B��Z���?m�����%���^f�'\��qRi��LYR-��ȼ&�m��w�c�ItR����'Uэ� �C���R����Wu�n5�^qO�����>|�,K۽������g�f�d����ͶpܪCLŷA���f��a�o�����)<K{�'h�8�k�A��=[~y�V����� +�繏�m�:�6������0�7*��Sm�����x�=uZ��-��9W����e��<�<�Bi�4}v�գ��J�vy��^Rɿ�F����Y�)����=��D��>�u�ǁ��WnZ<V؆��ۤ�*g��Z���Bi������/�,��@�CƗ��y����t˻N�-X�0m���nc�{g�#~�6��}I������|ʠ?����`<L�o����k������Q3*�ᑕ8}�1[����(f���-���b3K)0,����DGhqD�L����o�桦�f�_& ��:�h%��myn�ޮH�K+�1$�"9�@*h@�5)&�A!�*<��a\�.A�&]D��ǳ�v��h��JI<_��g����m��.���Dˋ�t�D%��C����:=L8ѡmF��	�id����P�+�4U:�n����o2�r�}�W�ᶽ	���cBJ!v{���V�67$���~��)�Y顄�i��܇U_�{�"�֟:M�W���zl��Ɍ!�#'��W}5"�ɑ�	SBە��뉠��r�2� �q�<�����'�(M�j�:���짒�U�ى����99�ghq�</��D���-�Y��+z'��C�"Y��s���L�h_�%�����o���)��� �f�t$RU�.<9�p�6�aa^��l�ԛ���EJ�e(�	,n>ZO	z�p�ì��G��_�� �V:����W�Wu*MC�'afda����"�ξ,H��t��RIiF�83��$����|�L��(��y�w�a�0m�������"��(����:|����)��>������:(
��7���@��*���@����6Hy�����R����4��@��-Q[6W��'7�O6��(,J�k#�o���%��Q�������H؎1��� R+�B�M���-�*����_�֓�Jd��)�v�)�SBR����3���� AQT����S}a�js/:7�����
�S��!=���%�.�(�ԋ��T�_jK*�3"-���"��=w֐��/�C�>ڌ�L���L1c�i�9N7�&���bլys� 
�T��n\�)���bi\7P�X)SC?m�j�{2�B�P� '�]Y& [~���UtF.��
��R|��ס�`w��c"�Oj�9��:��<�L��zj]onJ𙜅���yE�z�4��ޱ/J�Fm��A��Fگtf�*|�`�%F
8�:F���A H�Tk�[5����u�2�zis6E-�,q/A�9O)&r�B�0'տ=��v����V!�3�VA�R�{��5��z����>U��hC*
�q�e�݉r��$�e�Х�K*�����w\eB��d�Fm6[Y�G_�O��3�/���m�����6Cyi���IG��D���� ������]�\�����stY |G9�%zg����O�)�y�ι��ʥ�:�W��t�u�`V��񈞝ӵoNG�׎�}ۄ�Ўi�F�����hϩ�Gq;��I��L_�{#MS锫^F���6�"�3��Y���Zڙ%Hh�
�Bod���&� �zFe<�IGE`d�'�7�/����x:�����`,���Ꞥ��ɷ�|3N:vNE4���*�(!�RܗK,=�mdx���<�꿭v՟�Gr�>���#���9����8Q^6�I/Z
:l��;��'L;#4Ėf����iH;א��|ɾtM��0�bO")�����w��Kz�,��h\��_�DSaq��rp����]ߥԢ rP��)`� ���Ew`��S�I!|��&Ɛ�cj��L�#���