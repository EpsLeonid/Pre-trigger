XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Ұ)�L�8e#���m��L�M���k:��)>M4m��f��Ĝ�����W({]v��D�)�;���Fo,va��kb�H��А��W�;�/�'��;a`F����/��l#��tT��� b%�7h�1і޽]B>�'�NxtW�c�n��ߢ��C�e`/���WF6�A)e�J�=z>����R��?N$Ux�F�>a"��h+�#=v
�%���l��|�8�ǲ��[�fi�@�2x�V7���W��T疰ظ������}@��Q��$N�n��%�W����M�R�*�$ȯ�G1��jH.YN�N��^��N�ϊ��v�����T ]=�L�Jť�"�om�� ���z�@~-��hh#BKl~�ͨyí#�ny�Jd�[���ʚj8!���u���.N%U\���.o,m�1���ryT�K�~��)�+��=?�[�,�NB���PN0����|���;�b�5��*yF��`&M�?��G�Yn����eI0��I��]��ys6��v�Ř6�����{o;_F�$A��;|0;�.���8^�-`�+�_�.�Y�y���y�@��X*�-�����⧕�Pޤp1����;8"�-Ax�2�F���`[n��n�'�LM��c/-�C%����U[�����	H��5��7hR���þ�@����Lz����J�#%9��r�t�teğ�� Ɔ�b�R�ɤ3�"�Q�p�B[�p���n�҃��Q:MkV}�M�H�(�v��+(���c���XlxVHYEB    1111     710�Y��= r�����s�#\ͫ\�_,��nV��ف�*�R��霼��m�!�?�ǗrTv.�J�t�HwU�����WY�{�N>��4�f�����x�uezP�%�*_`�Mx�ٕ�E�7�͂pba��Ү$��$d���t�P�`n�>1��P1|-��ޚ��S��b,gz^Ak�C��b�i��8
ä�_-=���q|���i��υ�Jߍ�*k�[�)�h5�l��2C_NX+��l��|4��MO���ʂ��A)��Q<ẋ�\�·t?;o��r]�;}�y����I�Z�W�����#��h�<d�Y�FVe׋lOĽi���V~�p�xFQ���f�ɕ��:AdhA���`B]lfG�I��4��"�%�
�M�� 7�f@Ŭ�N��m�~�y�
7rg-]|�����3GG�&��O�
������;|a'�������c�+������.�b[��#VfS�� $�mc_\ �Ե��Cjv��u'VU����ЄK��aX�9��̶�p��@����Ŋ���>�`K��n�l��%�KS�8���q�V�UJ؝�w��}hS������{{��0��<(p1K�sS)O�)��V�m��Aqc m�^N�ឃ��?D�8�F��n�W<ک�Ə������Sx�D�E�px�ђp��1��k%$[G.��q�^��Bjg���>^��{�p$�|��Yu{���B�r�p_�B�[w�丮��i�rn'D�ְ��s��w撜�2EO��7���۽�o<2V���'�ō��'BG�:^0.��8>�����1���V*3Mq���
���c��D���_����A88�R(�@��G����H8>p�����_����A� K��^�Z�_�|�Z��O���,߈�RJb�f���~���P�^��!,ƅ��X�BD�V�m���	���lu��O���j*J������fUb�W���>��``^d�mn$Ad�ҽ�[�[���"LdP���a���r���<-���f�GM�6�!������z�K�R����0���o���%ns�5O�GN��bȥ�cU=�]������ԬxJ�0�5]FSV���k���p��*&O(Ԏτ���}���A�
8\�W���|d&��t'�9���vX�I�y�fGI�pT��kڈB3l;�xo�!Wm�G�$�l%�|������ �<�i.%�����|g�p�[�Y��@�ٰ���,=�lo&����)��	@w2�Fh�S �_��R�����ܯ7"o��!���gy3��t9���8n@n��<�E�#��tmLQ0@f���aQq���Gt� ��^�P����^B��'����6�� B��x���t@H��F,k�
U���C=}@�t~�vT�0�_���̹�G��?���ܥ��&Gr�zXE�z�!c����؈�A� ������
�D��nMd(�;۬1�v)�6I[�%v�E�.����:rp�G��Y����ჾ�[s+�|M����U}Yx7iFr�M��Y*�mIB ��T?i��1��YJ�+��T�iӁm�	���EF���V�3�ja��a��U�#�/�K�XkAzU����*Y��"�2Tʅ	�Wj��	-	v�G~���d�7l�J8�:I�<g52Yn��R$�P�%o� 	K��UR���Q��y}�ʰqQ���A���,:����U�y0���œg�3�#A�P(��P��SH�����?�:N���<�ͯ�ɴ<u!D9�)>廿S&u������	��