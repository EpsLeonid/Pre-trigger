XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D��^���Tį��&�S�g��e��:����H+��ID�R:���h��m�WUDG�j48��p���[�?��9�x�s�M�;�e��c�&(v�e���%����Y�cQ"�ӧo����&�R1�o�Yt��O`q紞݀AK�&����/��=�ų�:.k!����Y�h)�	&Q̅Z��Bw%t�;�4�6|�����5Y�dQ���h����A%V�GQ
a�Ї-�eS���	��?�0��rY��
J�5ك\�oL�U�dfh�d+����m�A�\)�$ c�U���Q+�3<�s��i3�s�o����q� i���t0�=��p��'洪�;�?��Tdx�~��Ւ�
�u�\�J0#�\l�����ٞ���M��A�����䲙�8���& �a(Zb_��M���p\QlS�4�<��C7�1.6r�(�Y�dQ뢚ICP�<p'�.�P�ݛ*�	��Kks�a<��n��}�/��qB�����KE����ϞD�(WO�6����>�Jh��V��[�=̩_�O�wz�4��B�'6S:��S�	���8����ҋ���ܯx=�V�4k~�Y���757�dϦ/��\PBB��]l��㦣�Wo���}�誴0�I[��$�ͣ��g�{^��7S�i����泵���x��ĝ
@�/�.���7����d�j�H���Є2
R� �S(��6Lu���||^�7�]���G���2�8<)yP�b'nSg�0��oB��	�ڗ|UXlxVHYEB    1eda     880E��i\B���cb�#��J��W�8�j
�u����5�rmj?�� ��*6s$c*��6�N��L�]O֣��hI���k$�"�M��ϔi<`�����xc�x�����ٛa�n}�X6� Y����p����;@1��sX�:���ih�/c���ޫ��M���d�+9��O��ٔ��n<�?m�څZU��n�\v��"}����:�Kj�WM�C��m�V��gӭw̠	�]����O�BKv{Jk�-����6�i���ޒ�g�-󰵰:��u��E �8����X}�a�Ӑo~�G��6��uw=��K��K���9I��\'V�X=�|ȇ�q�W��s���������}��a8��%�5����l�_���B��re52⍲ï���9�'�$0Ze�5+����D��+A}(��b���x[1�xB;&$�LcJF?5�dH�Nl�8�h֮v���Y,��"��Gٕ���jx�Rn�z��\�Thjo��Y�� 6�﫞���1(��j%sU��3���צ�P���nj�y�$!�e���];�iY��!���iw��Mfȧ#Ҥa1oH�~�xC6����/���a��b�떋M.0�Fq�Z�N�C�����ݩ�E����%�����Y�l�	g�o�\]v&6�x�����C҉�<E _�I�4�c=��Gu����Ar�O�y��]f��>�s�4�%���T�+2 �ޗ�@�	�um�a#`MI���E�?X�$����D<2ӷ���&�[+s�>	���q�<�6f,Y���i%HZ'��#E
���4d�g9�
���Vu����d�A;�
��gy���WA�4�w#�"Ź�u7B��Ε�WѷB�I�m�l$"E��gs�!_�9"�pI)�dT5W�x�.��7jl՝���݊�6�7ށ��|�z5Ʌ��>L�O����l��m溗�[v�̯xv` `a���~�:͟�נ�jn�ׇArzbe4#�=a��w8^����N�3�W,.>&��|&Ƹ�^�Bɲ�ϝ2�w�3J�[X�l�ۥ��E�-���!$�ԭ��;-��i�׫Ӱ̠d����,.wau��m�B�z{�؅��� �bp�:���3��n��}��C�6*�j5t�Ց��-;�6N+s���I��P�g���m���X�? �<(<�DK���&�����ƽN�b ���2�:�"@q�[�hp�L�F�D6	��3�V���cQ�+�{n�z.ו蠀	�O����%��u��:,�Hb	=��9 �S(@�������A��׺l&Ǿ�F���T�Z6 �-L�~�5/�S�m��&J�น���!��S��l��Џu&�Sê9� �k��\1u0�_�d��~�r�W���FI�Ӓ�N�uza�?��%�ޡ\X��I֖���s�G���޺/S�\E�9f�>���U���n��R9�N�T��E�_G���P�L�21MP1�8o�u̶D��@���f�ny5-�;�`9~;��7�Tv
���#�2���u@�^��:b��M�q�~�;��Ѯ�O�D���?�q��?� ��ZM��H���l�=b�k	�s6��M�e"���P�9TI�O�����Gm���j�yB'Q����|���(�Q��4<88�M�Ph�^���ڜ�䡌^����E��Ǖk��*��?���������6��q���.n|��P���]�)K�������n��-�<���j|\�|�D�	oU����4�cl�+:b�g�*�;V
Q�z���g��s�|�}Jq�I�+�%I�o
�V*���+�g�&:Gi��F+�Ć�%�� ψwק�ؠ�:#��t1���M�.
����1�i��?@*�Wꇆ�:r�h�hY֢�`�G;%A�c�y���/T��"L��)V�ל;��/\L=�k�gkiW-��$��TY��w�����j=���(�"���r��ѡ�5ފO�
�b�z�<��~~�)9}��m؛4��DM���E�f�[��7�3�#N.��~��2����S�w%�j��f;��[w����ir�d7����=�������g��^���;�[eڳ�Ȥ�,��������ZW��4*�Q�d��cS�M���K���t���qJ�D5c��C}.�������Ic��$�V�J�*�A���$ɽU 